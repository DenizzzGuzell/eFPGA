/*verilator tracing_on*/
//Example
//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Top-level Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed Aug 14 09:11:37 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype wire

// ----- Verilog module for fpga_top -----
module fpga_top(clk_i,
                Reset,
                prog_clk,
                IO_ISOL_N,
                gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN,
                gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT,
                gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR,
                ccff_head,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] clk_i;
//----- GLOBAL PORTS -----
input [0:0] Reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- GLOBAL PORTS -----
input [0:0] IO_ISOL_N;
//----- GPIN PORTS -----
input [0:143] gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN;
//----- GPOUT PORTS -----
output [0:143] gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT;
//----- GPOUT PORTS -----
output [0:143] gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR;
//----- INPUT PORTS -----
input [0:31] ccff_head;
//----- OUTPUT PORTS -----
output [0:31] ccff_tail;
/*verilator tracing_off*/
//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:0] direct_interc_0_out;
wire [0:0] direct_interc_100_out;
wire [0:0] direct_interc_101_out;
wire [0:0] direct_interc_102_out;
wire [0:0] direct_interc_103_out;
wire [0:0] direct_interc_104_out;
wire [0:0] direct_interc_105_out;
wire [0:0] direct_interc_106_out;
wire [0:0] direct_interc_107_out;
wire [0:0] direct_interc_108_out;
wire [0:0] direct_interc_109_out;
wire [0:0] direct_interc_10_out;
wire [0:0] direct_interc_110_out;
wire [0:0] direct_interc_111_out;
wire [0:0] direct_interc_112_out;
wire [0:0] direct_interc_113_out;
wire [0:0] direct_interc_114_out;
wire [0:0] direct_interc_115_out;
wire [0:0] direct_interc_116_out;
wire [0:0] direct_interc_117_out;
wire [0:0] direct_interc_118_out;
wire [0:0] direct_interc_119_out;
wire [0:0] direct_interc_11_out;
wire [0:0] direct_interc_120_out;
wire [0:0] direct_interc_121_out;
wire [0:0] direct_interc_122_out;
wire [0:0] direct_interc_123_out;
wire [0:0] direct_interc_124_out;
wire [0:0] direct_interc_125_out;
wire [0:0] direct_interc_126_out;
wire [0:0] direct_interc_127_out;
wire [0:0] direct_interc_128_out;
wire [0:0] direct_interc_129_out;
wire [0:0] direct_interc_12_out;
wire [0:0] direct_interc_130_out;
wire [0:0] direct_interc_131_out;
wire [0:0] direct_interc_132_out;
wire [0:0] direct_interc_133_out;
wire [0:0] direct_interc_134_out;
wire [0:0] direct_interc_135_out;
wire [0:0] direct_interc_136_out;
wire [0:0] direct_interc_137_out;
wire [0:0] direct_interc_138_out;
wire [0:0] direct_interc_139_out;
wire [0:0] direct_interc_13_out;
wire [0:0] direct_interc_140_out;
wire [0:0] direct_interc_141_out;
wire [0:0] direct_interc_142_out;
wire [0:0] direct_interc_143_out;
wire [0:0] direct_interc_144_out;
wire [0:0] direct_interc_145_out;
wire [0:0] direct_interc_146_out;
wire [0:0] direct_interc_147_out;
wire [0:0] direct_interc_148_out;
wire [0:0] direct_interc_149_out;
wire [0:0] direct_interc_14_out;
wire [0:0] direct_interc_150_out;
wire [0:0] direct_interc_151_out;
wire [0:0] direct_interc_152_out;
wire [0:0] direct_interc_153_out;
wire [0:0] direct_interc_154_out;
wire [0:0] direct_interc_155_out;
wire [0:0] direct_interc_156_out;
wire [0:0] direct_interc_157_out;
wire [0:0] direct_interc_158_out;
wire [0:0] direct_interc_159_out;
wire [0:0] direct_interc_15_out;
wire [0:0] direct_interc_160_out;
wire [0:0] direct_interc_161_out;
wire [0:0] direct_interc_162_out;
wire [0:0] direct_interc_163_out;
wire [0:0] direct_interc_164_out;
wire [0:0] direct_interc_165_out;
wire [0:0] direct_interc_166_out;
wire [0:0] direct_interc_167_out;
wire [0:0] direct_interc_168_out;
wire [0:0] direct_interc_169_out;
wire [0:0] direct_interc_16_out;
wire [0:0] direct_interc_170_out;
wire [0:0] direct_interc_171_out;
wire [0:0] direct_interc_172_out;
wire [0:0] direct_interc_173_out;
wire [0:0] direct_interc_174_out;
wire [0:0] direct_interc_175_out;
wire [0:0] direct_interc_176_out;
wire [0:0] direct_interc_177_out;
wire [0:0] direct_interc_178_out;
wire [0:0] direct_interc_179_out;
wire [0:0] direct_interc_17_out;
wire [0:0] direct_interc_180_out;
wire [0:0] direct_interc_181_out;
wire [0:0] direct_interc_182_out;
wire [0:0] direct_interc_183_out;
wire [0:0] direct_interc_184_out;
wire [0:0] direct_interc_185_out;
wire [0:0] direct_interc_186_out;
wire [0:0] direct_interc_187_out;
wire [0:0] direct_interc_188_out;
wire [0:0] direct_interc_189_out;
wire [0:0] direct_interc_18_out;
wire [0:0] direct_interc_190_out;
wire [0:0] direct_interc_191_out;
wire [0:0] direct_interc_192_out;
wire [0:0] direct_interc_193_out;
wire [0:0] direct_interc_194_out;
wire [0:0] direct_interc_195_out;
wire [0:0] direct_interc_196_out;
wire [0:0] direct_interc_197_out;
wire [0:0] direct_interc_19_out;
wire [0:0] direct_interc_1_out;
wire [0:0] direct_interc_20_out;
wire [0:0] direct_interc_21_out;
wire [0:0] direct_interc_22_out;
wire [0:0] direct_interc_23_out;
wire [0:0] direct_interc_24_out;
wire [0:0] direct_interc_25_out;
wire [0:0] direct_interc_26_out;
wire [0:0] direct_interc_27_out;
wire [0:0] direct_interc_28_out;
wire [0:0] direct_interc_29_out;
wire [0:0] direct_interc_2_out;
wire [0:0] direct_interc_30_out;
wire [0:0] direct_interc_31_out;
wire [0:0] direct_interc_32_out;
wire [0:0] direct_interc_33_out;
wire [0:0] direct_interc_34_out;
wire [0:0] direct_interc_35_out;
wire [0:0] direct_interc_36_out;
wire [0:0] direct_interc_37_out;
wire [0:0] direct_interc_38_out;
wire [0:0] direct_interc_39_out;
wire [0:0] direct_interc_3_out;
wire [0:0] direct_interc_40_out;
wire [0:0] direct_interc_41_out;
wire [0:0] direct_interc_42_out;
wire [0:0] direct_interc_43_out;
wire [0:0] direct_interc_44_out;
wire [0:0] direct_interc_45_out;
wire [0:0] direct_interc_46_out;
wire [0:0] direct_interc_47_out;
wire [0:0] direct_interc_48_out;
wire [0:0] direct_interc_49_out;
wire [0:0] direct_interc_4_out;
wire [0:0] direct_interc_50_out;
wire [0:0] direct_interc_51_out;
wire [0:0] direct_interc_52_out;
wire [0:0] direct_interc_53_out;
wire [0:0] direct_interc_54_out;
wire [0:0] direct_interc_55_out;
wire [0:0] direct_interc_56_out;
wire [0:0] direct_interc_57_out;
wire [0:0] direct_interc_58_out;
wire [0:0] direct_interc_59_out;
wire [0:0] direct_interc_5_out;
wire [0:0] direct_interc_60_out;
wire [0:0] direct_interc_61_out;
wire [0:0] direct_interc_62_out;
wire [0:0] direct_interc_63_out;
wire [0:0] direct_interc_64_out;
wire [0:0] direct_interc_65_out;
wire [0:0] direct_interc_66_out;
wire [0:0] direct_interc_67_out;
wire [0:0] direct_interc_68_out;
wire [0:0] direct_interc_69_out;
wire [0:0] direct_interc_6_out;
wire [0:0] direct_interc_70_out;
wire [0:0] direct_interc_71_out;
wire [0:0] direct_interc_72_out;
wire [0:0] direct_interc_73_out;
wire [0:0] direct_interc_74_out;
wire [0:0] direct_interc_75_out;
wire [0:0] direct_interc_76_out;
wire [0:0] direct_interc_77_out;
wire [0:0] direct_interc_78_out;
wire [0:0] direct_interc_79_out;
wire [0:0] direct_interc_7_out;
wire [0:0] direct_interc_80_out;
wire [0:0] direct_interc_81_out;
wire [0:0] direct_interc_82_out;
wire [0:0] direct_interc_83_out;
wire [0:0] direct_interc_84_out;
wire [0:0] direct_interc_85_out;
wire [0:0] direct_interc_86_out;
wire [0:0] direct_interc_87_out;
wire [0:0] direct_interc_88_out;
wire [0:0] direct_interc_89_out;
wire [0:0] direct_interc_8_out;
wire [0:0] direct_interc_90_out;
wire [0:0] direct_interc_91_out;
wire [0:0] direct_interc_92_out;
wire [0:0] direct_interc_93_out;
wire [0:0] direct_interc_94_out;
wire [0:0] direct_interc_95_out;
wire [0:0] direct_interc_96_out;
wire [0:0] direct_interc_97_out;
wire [0:0] direct_interc_98_out;
wire [0:0] direct_interc_99_out;
wire [0:0] direct_interc_9_out;
wire [0:64] tile_0__10__0_cby_0__10__chany_top_out;
wire [0:0] tile_0__10__0_ccff_tail;
wire [0:0] tile_0__10__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__10__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__10__0_sb_0__9__chanx_right_out;
wire [0:64] tile_0__10__0_sb_0__9__chany_bottom_out;
wire [0:64] tile_0__11__0_cby_0__11__chany_top_out;
wire [0:0] tile_0__11__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__11__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__11__0_sb_0__10__chanx_right_out;
wire [0:64] tile_0__11__0_sb_0__10__chany_bottom_out;
wire [0:64] tile_0__19__0_sb_0__18__chanx_right_out;
wire [0:64] tile_0__19__0_sb_0__18__chany_bottom_out;
wire [0:64] tile_0__1__0_cby_0__1__chany_top_out;
wire [0:0] tile_0__1__0_ccff_tail;
wire [0:0] tile_0__1__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__1__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__1__0_sb_0__0__chanx_right_out;
wire [0:64] tile_0__2__0_cby_0__2__chany_top_out;
wire [0:0] tile_0__2__0_ccff_tail;
wire [0:0] tile_0__2__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__2__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__2__0_sb_0__1__chanx_right_out;
wire [0:64] tile_0__2__0_sb_0__1__chany_bottom_out;
wire [0:64] tile_0__2__10_cby_0__2__chany_top_out;
wire [0:0] tile_0__2__10_ccff_tail;
wire [0:0] tile_0__2__10_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__2__10_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__2__10_sb_0__1__chanx_right_out;
wire [0:64] tile_0__2__10_sb_0__1__chany_bottom_out;
wire [0:64] tile_0__2__1_cby_0__2__chany_top_out;
wire [0:0] tile_0__2__1_ccff_tail;
wire [0:0] tile_0__2__1_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__2__1_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__2__1_sb_0__1__chanx_right_out;
wire [0:64] tile_0__2__1_sb_0__1__chany_bottom_out;
wire [0:64] tile_0__2__2_cby_0__2__chany_top_out;
wire [0:0] tile_0__2__2_ccff_tail;
wire [0:0] tile_0__2__2_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__2__2_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__2__2_sb_0__1__chanx_right_out;
wire [0:64] tile_0__2__2_sb_0__1__chany_bottom_out;
wire [0:64] tile_0__2__3_cby_0__2__chany_top_out;
wire [0:0] tile_0__2__3_ccff_tail;
wire [0:0] tile_0__2__3_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__2__3_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__2__3_sb_0__1__chanx_right_out;
wire [0:64] tile_0__2__3_sb_0__1__chany_bottom_out;
wire [0:64] tile_0__2__4_cby_0__2__chany_top_out;
wire [0:0] tile_0__2__4_ccff_tail;
wire [0:0] tile_0__2__4_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__2__4_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__2__4_sb_0__1__chanx_right_out;
wire [0:64] tile_0__2__4_sb_0__1__chany_bottom_out;
wire [0:64] tile_0__2__5_cby_0__2__chany_top_out;
wire [0:0] tile_0__2__5_ccff_tail;
wire [0:0] tile_0__2__5_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__2__5_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__2__5_sb_0__1__chanx_right_out;
wire [0:64] tile_0__2__5_sb_0__1__chany_bottom_out;
wire [0:64] tile_0__2__6_cby_0__2__chany_top_out;
wire [0:0] tile_0__2__6_ccff_tail;
wire [0:0] tile_0__2__6_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__2__6_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__2__6_sb_0__1__chanx_right_out;
wire [0:64] tile_0__2__6_sb_0__1__chany_bottom_out;
wire [0:64] tile_0__2__7_cby_0__2__chany_top_out;
wire [0:0] tile_0__2__7_ccff_tail;
wire [0:0] tile_0__2__7_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__2__7_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__2__7_sb_0__1__chanx_right_out;
wire [0:64] tile_0__2__7_sb_0__1__chany_bottom_out;
wire [0:64] tile_0__2__8_cby_0__2__chany_top_out;
wire [0:0] tile_0__2__8_ccff_tail;
wire [0:0] tile_0__2__8_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__2__8_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__2__8_sb_0__1__chanx_right_out;
wire [0:64] tile_0__2__8_sb_0__1__chany_bottom_out;
wire [0:64] tile_0__2__9_cby_0__2__chany_top_out;
wire [0:0] tile_0__2__9_ccff_tail;
wire [0:0] tile_0__2__9_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__2__9_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__2__9_sb_0__1__chanx_right_out;
wire [0:64] tile_0__2__9_sb_0__1__chany_bottom_out;
wire [0:64] tile_0__5__0_cby_0__5__chany_top_out;
wire [0:0] tile_0__5__0_ccff_tail;
wire [0:0] tile_0__5__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__5__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__5__0_sb_0__4__chanx_right_out;
wire [0:64] tile_0__5__0_sb_0__4__chany_bottom_out;
wire [0:64] tile_0__5__1_cby_0__5__chany_top_out;
wire [0:0] tile_0__5__1_ccff_tail;
wire [0:0] tile_0__5__1_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__5__1_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__5__1_sb_0__4__chanx_right_out;
wire [0:64] tile_0__5__1_sb_0__4__chany_bottom_out;
wire [0:64] tile_0__6__0_cby_0__6__chany_top_out;
wire [0:0] tile_0__6__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__6__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__6__0_sb_0__5__chanx_right_out;
wire [0:64] tile_0__6__0_sb_0__5__chany_bottom_out;
wire [0:64] tile_0__6__1_cby_0__6__chany_top_out;
wire [0:0] tile_0__6__1_ccff_tail;
wire [0:0] tile_0__6__1_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__6__1_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__6__1_sb_0__5__chanx_right_out;
wire [0:64] tile_0__6__1_sb_0__5__chany_bottom_out;
wire [0:0] tile_10__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_10__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_10__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_10__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_10__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_10__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_10__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_10__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_11__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_11__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_11__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_11__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_11__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_11__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_11__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_11__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_12__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_12__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_12__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_12__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_12__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_12__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_12__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_12__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_13__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_13__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_13__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_13__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_13__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_13__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_13__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_13__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_14__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_14__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_14__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_14__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_14__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_14__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_14__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_14__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_15__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_15__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_15__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_15__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_15__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_15__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_15__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_15__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_16__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_16__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_16__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_16__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_16__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_16__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_16__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_16__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_17__10__0_cbx_17__9__chanx_left_out;
wire [0:0] tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_17__10__0_cby_18__10__chany_top_out;
wire [0:0] tile_17__10__0_cby_18__10__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_17__10__0_cby_18__10__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_17__10__0_ccff_tail;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_;
wire [0:64] tile_17__10__0_sb_17__9__chany_bottom_out;
wire [0:64] tile_17__10__0_sb_18__9__chany_bottom_out;
wire [0:0] tile_17__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_17__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_17__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_17__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_17__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_17__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_17__5__0_cbx_17__4__chanx_left_out;
wire [0:0] tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_17__5__0_cby_18__5__chany_top_out;
wire [0:0] tile_17__5__0_cby_18__5__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_17__5__0_cby_18__5__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_17__5__0_ccff_tail;
wire [0:0] tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_17__5__0_sb_17__4__chany_bottom_out;
wire [0:64] tile_17__5__0_sb_18__4__chany_bottom_out;
wire [0:0] tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_17__5__1_cbx_17__4__chanx_left_out;
wire [0:0] tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_17__5__1_cby_18__5__chany_top_out;
wire [0:0] tile_17__5__1_cby_18__5__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_17__5__1_cby_18__5__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_17__5__1_ccff_tail;
wire [0:0] tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_17__5__1_sb_17__4__chany_bottom_out;
wire [0:64] tile_17__5__1_sb_18__4__chany_bottom_out;
wire [0:0] tile_17__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_17__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_18__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_18__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_18__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_18__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_18__19__0_cbx_18__18__chanx_left_out;
wire [0:0] tile_18__19__0_ccff_tail;
wire [0:0] tile_18__19__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_18__19__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_18__19__0_sb_18__18__chany_bottom_out;
wire [0:0] tile_18__1__0_cbx_18__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_18__1__0_cbx_18__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_18__1__0_cbx_18__0__chanx_left_out;
wire [0:64] tile_18__1__0_cby_18__1__chany_top_out;
wire [0:0] tile_18__1__0_cby_18__1__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_18__1__0_cby_18__1__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_18__1__0_ccff_tail;
wire [0:0] tile_18__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_18__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_18__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_18__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_18__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_18__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_18__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_18__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_18__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_18__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] tile_18__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_18__2__0_cbx_18__1__chanx_left_out;
wire [0:64] tile_18__2__0_cby_18__2__chany_top_out;
wire [0:0] tile_18__2__0_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_18__2__0_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_18__2__0_ccff_tail;
wire [0:0] tile_18__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_18__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_18__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_18__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_18__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_18__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_18__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_18__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_18__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_18__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_18__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_18__2__0_sb_18__1__chany_bottom_out;
wire [0:0] tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_18__2__10_cbx_18__1__chanx_left_out;
wire [0:64] tile_18__2__10_cby_18__2__chany_top_out;
wire [0:0] tile_18__2__10_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_18__2__10_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_18__2__10_ccff_tail;
wire [0:0] tile_18__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_18__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_18__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_18__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_18__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_18__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_18__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_18__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_18__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_18__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_18__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_18__2__10_sb_18__1__chany_bottom_out;
wire [0:0] tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_18__2__1_cbx_18__1__chanx_left_out;
wire [0:64] tile_18__2__1_cby_18__2__chany_top_out;
wire [0:0] tile_18__2__1_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_18__2__1_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_18__2__1_ccff_tail;
wire [0:0] tile_18__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_18__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_18__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_18__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_18__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_18__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_18__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_18__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_18__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_18__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_18__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_18__2__1_sb_18__1__chany_bottom_out;
wire [0:0] tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_18__2__2_cbx_18__1__chanx_left_out;
wire [0:64] tile_18__2__2_cby_18__2__chany_top_out;
wire [0:0] tile_18__2__2_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_18__2__2_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_18__2__2_ccff_tail;
wire [0:0] tile_18__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_18__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_18__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_18__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_18__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_18__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_18__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_18__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_18__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_18__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_18__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_18__2__2_sb_18__1__chany_bottom_out;
wire [0:0] tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_18__2__3_cbx_18__1__chanx_left_out;
wire [0:64] tile_18__2__3_cby_18__2__chany_top_out;
wire [0:0] tile_18__2__3_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_18__2__3_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_18__2__3_ccff_tail;
wire [0:0] tile_18__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_18__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_18__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_18__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_18__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_18__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_18__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_18__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_18__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_18__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_18__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_18__2__3_sb_18__1__chany_bottom_out;
wire [0:0] tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_18__2__4_cbx_18__1__chanx_left_out;
wire [0:64] tile_18__2__4_cby_18__2__chany_top_out;
wire [0:0] tile_18__2__4_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_18__2__4_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_18__2__4_ccff_tail;
wire [0:0] tile_18__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_18__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_18__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_18__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_18__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_18__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_18__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_18__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_18__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_18__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_18__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_18__2__4_sb_18__1__chany_bottom_out;
wire [0:0] tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_18__2__5_cbx_18__1__chanx_left_out;
wire [0:64] tile_18__2__5_cby_18__2__chany_top_out;
wire [0:0] tile_18__2__5_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_18__2__5_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_18__2__5_ccff_tail;
wire [0:0] tile_18__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_18__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_18__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_18__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_18__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_18__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_18__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_18__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_18__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_18__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_18__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_18__2__5_sb_18__1__chany_bottom_out;
wire [0:0] tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_18__2__6_cbx_18__1__chanx_left_out;
wire [0:64] tile_18__2__6_cby_18__2__chany_top_out;
wire [0:0] tile_18__2__6_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_18__2__6_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_18__2__6_ccff_tail;
wire [0:0] tile_18__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_18__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_18__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_18__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_18__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_18__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_18__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_18__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_18__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_18__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_18__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_18__2__6_sb_18__1__chany_bottom_out;
wire [0:0] tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_18__2__7_cbx_18__1__chanx_left_out;
wire [0:64] tile_18__2__7_cby_18__2__chany_top_out;
wire [0:0] tile_18__2__7_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_18__2__7_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_18__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_18__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_18__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_18__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_18__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_18__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_18__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_18__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_18__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_18__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_18__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_18__2__7_sb_18__1__chany_bottom_out;
wire [0:0] tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_18__2__8_cbx_18__1__chanx_left_out;
wire [0:64] tile_18__2__8_cby_18__2__chany_top_out;
wire [0:0] tile_18__2__8_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_18__2__8_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_18__2__8_ccff_tail;
wire [0:0] tile_18__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_18__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_18__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_18__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_18__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_18__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_18__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_18__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_18__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_18__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_18__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_18__2__8_sb_18__1__chany_bottom_out;
wire [0:0] tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_18__2__9_cbx_18__1__chanx_left_out;
wire [0:64] tile_18__2__9_cby_18__2__chany_top_out;
wire [0:0] tile_18__2__9_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_18__2__9_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_18__2__9_ccff_tail;
wire [0:0] tile_18__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_18__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_18__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_18__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_18__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_18__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_18__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_18__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_18__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_18__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_18__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_18__2__9_sb_18__1__chany_bottom_out;
wire [0:0] tile_18__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:64] tile_18__6__0_cbx_18__5__chanx_left_out;
wire [0:64] tile_18__6__0_cby_18__6__chany_top_out;
wire [0:0] tile_18__6__0_cby_18__6__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_18__6__0_cby_18__6__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_18__6__0_ccff_tail;
wire [0:0] tile_18__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_18__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_18__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_18__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_18__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_18__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_18__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_18__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_18__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_18__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_18__6__0_sb_18__5__chany_bottom_out;
wire [0:64] tile_18__6__1_cbx_18__5__chanx_left_out;
wire [0:64] tile_18__6__1_cby_18__6__chany_top_out;
wire [0:0] tile_18__6__1_cby_18__6__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_18__6__1_cby_18__6__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_18__6__1_ccff_tail;
wire [0:0] tile_18__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_18__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_18__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_18__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_18__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_18__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_18__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_18__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_18__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_18__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_18__6__1_sb_18__5__chany_bottom_out;
wire [0:64] tile_18__6__2_cbx_18__5__chanx_left_out;
wire [0:64] tile_18__6__2_cby_18__6__chany_top_out;
wire [0:0] tile_18__6__2_cby_18__6__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_18__6__2_cby_18__6__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_18__6__2_ccff_tail;
wire [0:0] tile_18__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_18__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_18__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_18__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_18__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_18__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_18__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_18__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_18__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_18__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_18__6__2_sb_18__5__chany_bottom_out;
wire [0:0] tile_18__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_18__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_19__1__0_ccff_tail;
wire [0:0] tile_19__1__0_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_19__1__0_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_19__1__10_ccff_tail;
wire [0:0] tile_19__1__10_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_19__1__10_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_19__1__11_ccff_tail;
wire [0:0] tile_19__1__11_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_19__1__11_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_19__1__12_ccff_tail;
wire [0:0] tile_19__1__12_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_19__1__12_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_19__1__13_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_19__1__13_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_19__1__14_ccff_tail;
wire [0:0] tile_19__1__14_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_19__1__14_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_19__1__15_ccff_tail;
wire [0:0] tile_19__1__15_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_19__1__15_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_19__1__16_ccff_tail;
wire [0:0] tile_19__1__16_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_19__1__16_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_19__1__17_ccff_tail;
wire [0:0] tile_19__1__17_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_19__1__17_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_19__1__1_ccff_tail;
wire [0:0] tile_19__1__1_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_19__1__1_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_19__1__2_ccff_tail;
wire [0:0] tile_19__1__2_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_19__1__2_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_19__1__3_ccff_tail;
wire [0:0] tile_19__1__3_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_19__1__3_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_19__1__4_ccff_tail;
wire [0:0] tile_19__1__4_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_19__1__4_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_19__1__5_ccff_tail;
wire [0:0] tile_19__1__5_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_19__1__5_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_19__1__6_ccff_tail;
wire [0:0] tile_19__1__6_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_19__1__6_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_19__1__7_ccff_tail;
wire [0:0] tile_19__1__7_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_19__1__7_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_19__1__8_ccff_tail;
wire [0:0] tile_19__1__8_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_19__1__8_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_19__1__9_ccff_tail;
wire [0:0] tile_19__1__9_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_19__1__9_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__0_ccff_tail;
wire [0:0] tile_1__0__0_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__0_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__10_ccff_tail;
wire [0:0] tile_1__0__10_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__10_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__11_ccff_tail;
wire [0:0] tile_1__0__11_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__11_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__12_ccff_tail;
wire [0:0] tile_1__0__12_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__12_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__13_ccff_tail;
wire [0:0] tile_1__0__13_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__13_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__14_ccff_tail;
wire [0:0] tile_1__0__14_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__14_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__15_ccff_tail;
wire [0:0] tile_1__0__15_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__15_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__16_ccff_tail;
wire [0:0] tile_1__0__16_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__16_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__17_ccff_tail;
wire [0:0] tile_1__0__17_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__17_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__1_ccff_tail;
wire [0:0] tile_1__0__1_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__1_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__2_ccff_tail;
wire [0:0] tile_1__0__2_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__2_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__3_ccff_tail;
wire [0:0] tile_1__0__3_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__3_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__4_ccff_tail;
wire [0:0] tile_1__0__4_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__4_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__5_ccff_tail;
wire [0:0] tile_1__0__5_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__5_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__6_ccff_tail;
wire [0:0] tile_1__0__6_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__6_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__7_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__7_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__8_ccff_tail;
wire [0:0] tile_1__0__8_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__8_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__9_ccff_tail;
wire [0:0] tile_1__0__9_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__9_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__10__0_cbx_1__9__chanx_left_out;
wire [0:0] tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__10__0_cby_2__10__chany_top_out;
wire [0:0] tile_1__10__0_ccff_tail;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_;
wire [0:64] tile_1__10__0_sb_1__9__chany_bottom_out;
wire [0:64] tile_1__10__0_sb_2__9__chanx_right_out;
wire [0:64] tile_1__10__0_sb_2__9__chany_bottom_out;
wire [0:0] tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__10__1_cbx_1__9__chanx_left_out;
wire [0:0] tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__10__1_cby_2__10__chany_top_out;
wire [0:0] tile_1__10__1_ccff_tail;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_;
wire [0:64] tile_1__10__1_sb_1__9__chany_bottom_out;
wire [0:64] tile_1__10__1_sb_2__9__chanx_right_out;
wire [0:64] tile_1__10__1_sb_2__9__chany_bottom_out;
wire [0:0] tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__10__2_cbx_1__9__chanx_left_out;
wire [0:0] tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__10__2_cby_2__10__chany_top_out;
wire [0:0] tile_1__10__2_ccff_tail;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_;
wire [0:64] tile_1__10__2_sb_1__9__chany_bottom_out;
wire [0:64] tile_1__10__2_sb_2__9__chanx_right_out;
wire [0:64] tile_1__10__2_sb_2__9__chany_bottom_out;
wire [0:0] tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__10__3_cbx_1__9__chanx_left_out;
wire [0:0] tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__10__3_cby_2__10__chany_top_out;
wire [0:0] tile_1__10__3_ccff_tail;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_;
wire [0:64] tile_1__10__3_sb_1__9__chany_bottom_out;
wire [0:64] tile_1__10__3_sb_2__9__chanx_right_out;
wire [0:64] tile_1__10__3_sb_2__9__chany_bottom_out;
wire [0:0] tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__10__4_cbx_1__9__chanx_left_out;
wire [0:0] tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__10__4_cby_2__10__chany_top_out;
wire [0:0] tile_1__10__4_ccff_tail;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_;
wire [0:64] tile_1__10__4_sb_1__9__chany_bottom_out;
wire [0:64] tile_1__10__4_sb_2__9__chanx_right_out;
wire [0:64] tile_1__10__4_sb_2__9__chany_bottom_out;
wire [0:0] tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__10__5_cbx_1__9__chanx_left_out;
wire [0:0] tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__10__5_cby_2__10__chany_top_out;
wire [0:0] tile_1__10__5_ccff_tail;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_;
wire [0:64] tile_1__10__5_sb_1__9__chany_bottom_out;
wire [0:64] tile_1__10__5_sb_2__9__chanx_right_out;
wire [0:64] tile_1__10__5_sb_2__9__chany_bottom_out;
wire [0:0] tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__10__6_cbx_1__9__chanx_left_out;
wire [0:0] tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__10__6_cby_2__10__chany_top_out;
wire [0:0] tile_1__10__6_ccff_tail;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_;
wire [0:64] tile_1__10__6_sb_1__9__chany_bottom_out;
wire [0:64] tile_1__10__6_sb_2__9__chanx_right_out;
wire [0:64] tile_1__10__6_sb_2__9__chany_bottom_out;
wire [0:0] tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__10__7_cbx_1__9__chanx_left_out;
wire [0:0] tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__10__7_cby_2__10__chany_top_out;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_;
wire [0:64] tile_1__10__7_sb_1__9__chany_bottom_out;
wire [0:64] tile_1__10__7_sb_2__9__chanx_right_out;
wire [0:64] tile_1__10__7_sb_2__9__chany_bottom_out;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_;
wire [0:0] tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_;
wire [0:64] tile_1__11__0_cbx_1__10__chanx_left_out;
wire [0:64] tile_1__11__0_cby_1__11__chany_top_out;
wire [0:0] tile_1__11__0_ccff_tail;
wire [0:0] tile_1__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__11__0_sb_1__10__chanx_right_out;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_;
wire [0:0] tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_;
wire [0:64] tile_1__11__1_cbx_1__10__chanx_left_out;
wire [0:64] tile_1__11__1_cby_1__11__chany_top_out;
wire [0:0] tile_1__11__1_ccff_tail;
wire [0:0] tile_1__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__11__1_sb_1__10__chanx_right_out;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_;
wire [0:0] tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_;
wire [0:64] tile_1__11__2_cbx_1__10__chanx_left_out;
wire [0:64] tile_1__11__2_cby_1__11__chany_top_out;
wire [0:0] tile_1__11__2_ccff_tail;
wire [0:0] tile_1__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__11__2_sb_1__10__chanx_right_out;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_;
wire [0:0] tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_;
wire [0:64] tile_1__11__3_cbx_1__10__chanx_left_out;
wire [0:64] tile_1__11__3_cby_1__11__chany_top_out;
wire [0:0] tile_1__11__3_ccff_tail;
wire [0:0] tile_1__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__11__3_sb_1__10__chanx_right_out;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_;
wire [0:0] tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_;
wire [0:64] tile_1__11__4_cbx_1__10__chanx_left_out;
wire [0:64] tile_1__11__4_cby_1__11__chany_top_out;
wire [0:0] tile_1__11__4_ccff_tail;
wire [0:0] tile_1__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__11__4_sb_1__10__chanx_right_out;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_;
wire [0:0] tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_;
wire [0:64] tile_1__11__5_cbx_1__10__chanx_left_out;
wire [0:64] tile_1__11__5_cby_1__11__chany_top_out;
wire [0:0] tile_1__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__11__5_sb_1__10__chanx_right_out;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_;
wire [0:0] tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_;
wire [0:64] tile_1__11__6_cbx_1__10__chanx_left_out;
wire [0:64] tile_1__11__6_cby_1__11__chany_top_out;
wire [0:0] tile_1__11__6_ccff_tail;
wire [0:0] tile_1__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__11__6_sb_1__10__chanx_right_out;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_;
wire [0:0] tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_;
wire [0:64] tile_1__11__7_cbx_1__10__chanx_left_out;
wire [0:64] tile_1__11__7_cby_1__11__chany_top_out;
wire [0:0] tile_1__11__7_ccff_tail;
wire [0:0] tile_1__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__11__7_sb_1__10__chanx_right_out;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_;
wire [0:0] tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_;
wire [0:64] tile_1__11__8_cbx_1__10__chanx_left_out;
wire [0:64] tile_1__11__8_cby_1__11__chany_top_out;
wire [0:0] tile_1__11__8_ccff_tail;
wire [0:0] tile_1__11__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__11__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__11__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__11__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__11__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__11__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__11__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__11__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__11__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__11__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__11__8_sb_1__10__chanx_right_out;
wire [0:0] tile_1__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_1__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__19__0_cbx_1__18__chanx_left_out;
wire [0:0] tile_1__19__0_ccff_tail;
wire [0:0] tile_1__19__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__19__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_1__19__0_sb_1__18__chanx_right_out;
wire [0:64] tile_1__19__0_sb_1__18__chany_bottom_out;
wire [0:0] tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__19__10_cbx_1__18__chanx_left_out;
wire [0:0] tile_1__19__10_ccff_tail;
wire [0:0] tile_1__19__10_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__19__10_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_1__19__10_sb_1__18__chanx_right_out;
wire [0:64] tile_1__19__10_sb_1__18__chany_bottom_out;
wire [0:0] tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__19__11_cbx_1__18__chanx_left_out;
wire [0:0] tile_1__19__11_ccff_tail;
wire [0:0] tile_1__19__11_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__19__11_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_1__19__11_sb_1__18__chanx_right_out;
wire [0:64] tile_1__19__11_sb_1__18__chany_bottom_out;
wire [0:0] tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__19__12_cbx_1__18__chanx_left_out;
wire [0:0] tile_1__19__12_ccff_tail;
wire [0:0] tile_1__19__12_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__19__12_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_1__19__12_sb_1__18__chanx_right_out;
wire [0:64] tile_1__19__12_sb_1__18__chany_bottom_out;
wire [0:0] tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__19__13_cbx_1__18__chanx_left_out;
wire [0:0] tile_1__19__13_ccff_tail;
wire [0:0] tile_1__19__13_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__19__13_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_1__19__13_sb_1__18__chanx_right_out;
wire [0:64] tile_1__19__13_sb_1__18__chany_bottom_out;
wire [0:0] tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__19__14_cbx_1__18__chanx_left_out;
wire [0:0] tile_1__19__14_ccff_tail;
wire [0:0] tile_1__19__14_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__19__14_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_1__19__14_sb_1__18__chanx_right_out;
wire [0:64] tile_1__19__14_sb_1__18__chany_bottom_out;
wire [0:0] tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__19__15_cbx_1__18__chanx_left_out;
wire [0:0] tile_1__19__15_ccff_tail;
wire [0:0] tile_1__19__15_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__19__15_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_1__19__15_sb_1__18__chanx_right_out;
wire [0:64] tile_1__19__15_sb_1__18__chany_bottom_out;
wire [0:0] tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__19__16_cbx_1__18__chanx_left_out;
wire [0:0] tile_1__19__16_ccff_tail;
wire [0:0] tile_1__19__16_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__19__16_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_1__19__16_sb_1__18__chanx_right_out;
wire [0:64] tile_1__19__16_sb_1__18__chany_bottom_out;
wire [0:0] tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__19__1_cbx_1__18__chanx_left_out;
wire [0:0] tile_1__19__1_ccff_tail;
wire [0:0] tile_1__19__1_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__19__1_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_1__19__1_sb_1__18__chanx_right_out;
wire [0:64] tile_1__19__1_sb_1__18__chany_bottom_out;
wire [0:0] tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__19__2_cbx_1__18__chanx_left_out;
wire [0:0] tile_1__19__2_ccff_tail;
wire [0:0] tile_1__19__2_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__19__2_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_1__19__2_sb_1__18__chanx_right_out;
wire [0:64] tile_1__19__2_sb_1__18__chany_bottom_out;
wire [0:0] tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__19__3_cbx_1__18__chanx_left_out;
wire [0:0] tile_1__19__3_ccff_tail;
wire [0:0] tile_1__19__3_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__19__3_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_1__19__3_sb_1__18__chanx_right_out;
wire [0:64] tile_1__19__3_sb_1__18__chany_bottom_out;
wire [0:0] tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__19__4_cbx_1__18__chanx_left_out;
wire [0:0] tile_1__19__4_ccff_tail;
wire [0:0] tile_1__19__4_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__19__4_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_1__19__4_sb_1__18__chanx_right_out;
wire [0:64] tile_1__19__4_sb_1__18__chany_bottom_out;
wire [0:0] tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__19__5_cbx_1__18__chanx_left_out;
wire [0:0] tile_1__19__5_ccff_tail;
wire [0:0] tile_1__19__5_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__19__5_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_1__19__5_sb_1__18__chanx_right_out;
wire [0:64] tile_1__19__5_sb_1__18__chany_bottom_out;
wire [0:0] tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__19__6_cbx_1__18__chanx_left_out;
wire [0:0] tile_1__19__6_ccff_tail;
wire [0:0] tile_1__19__6_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__19__6_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_1__19__6_sb_1__18__chanx_right_out;
wire [0:64] tile_1__19__6_sb_1__18__chany_bottom_out;
wire [0:0] tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__19__7_cbx_1__18__chanx_left_out;
wire [0:0] tile_1__19__7_ccff_tail;
wire [0:0] tile_1__19__7_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__19__7_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_1__19__7_sb_1__18__chanx_right_out;
wire [0:64] tile_1__19__7_sb_1__18__chany_bottom_out;
wire [0:0] tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__19__8_cbx_1__18__chanx_left_out;
wire [0:0] tile_1__19__8_ccff_tail;
wire [0:0] tile_1__19__8_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__19__8_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_1__19__8_sb_1__18__chanx_right_out;
wire [0:64] tile_1__19__8_sb_1__18__chany_bottom_out;
wire [0:0] tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__19__9_cbx_1__18__chanx_left_out;
wire [0:0] tile_1__19__9_ccff_tail;
wire [0:0] tile_1__19__9_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__19__9_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_1__19__9_sb_1__18__chanx_right_out;
wire [0:64] tile_1__19__9_sb_1__18__chany_bottom_out;
wire [0:0] tile_1__1__0_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_1__1__0_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_1__1__0_cbx_1__0__chanx_left_out;
wire [0:64] tile_1__1__0_cby_1__1__chany_top_out;
wire [0:0] tile_1__1__0_ccff_tail;
wire [0:0] tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__1__0_sb_1__0__chanx_right_out;
wire [0:0] tile_1__1__10_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_1__1__10_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_1__1__10_cbx_1__0__chanx_left_out;
wire [0:64] tile_1__1__10_cby_1__1__chany_top_out;
wire [0:0] tile_1__1__10_ccff_tail;
wire [0:0] tile_1__1__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__1__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__1__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__1__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__1__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__1__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__1__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__1__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__1__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__1__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__1__10_sb_1__0__chanx_right_out;
wire [0:0] tile_1__1__11_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_1__1__11_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_1__1__11_cbx_1__0__chanx_left_out;
wire [0:64] tile_1__1__11_cby_1__1__chany_top_out;
wire [0:0] tile_1__1__11_ccff_tail;
wire [0:0] tile_1__1__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__1__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__1__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__1__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__1__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__1__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__1__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__1__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__1__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__1__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__1__11_sb_1__0__chanx_right_out;
wire [0:0] tile_1__1__12_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_1__1__12_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_1__1__12_cbx_1__0__chanx_left_out;
wire [0:64] tile_1__1__12_cby_1__1__chany_top_out;
wire [0:0] tile_1__1__12_ccff_tail;
wire [0:0] tile_1__1__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__1__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__1__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__1__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__1__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__1__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__1__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__1__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__1__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__1__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__1__12_sb_1__0__chanx_right_out;
wire [0:0] tile_1__1__13_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_1__1__13_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_1__1__13_cbx_1__0__chanx_left_out;
wire [0:64] tile_1__1__13_cby_1__1__chany_top_out;
wire [0:0] tile_1__1__13_ccff_tail;
wire [0:0] tile_1__1__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__1__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__1__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__1__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__1__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__1__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__1__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__1__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__1__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__1__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__1__13_sb_1__0__chanx_right_out;
wire [0:0] tile_1__1__14_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_1__1__14_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_1__1__14_cbx_1__0__chanx_left_out;
wire [0:64] tile_1__1__14_cby_1__1__chany_top_out;
wire [0:0] tile_1__1__14_ccff_tail;
wire [0:0] tile_1__1__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__1__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__1__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__1__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__1__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__1__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__1__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__1__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__1__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__1__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__1__14_sb_1__0__chanx_right_out;
wire [0:0] tile_1__1__15_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_1__1__15_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_1__1__15_cbx_1__0__chanx_left_out;
wire [0:64] tile_1__1__15_cby_1__1__chany_top_out;
wire [0:0] tile_1__1__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__1__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__1__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__1__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__1__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__1__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__1__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__1__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__1__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__1__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__1__15_sb_1__0__chanx_right_out;
wire [0:0] tile_1__1__16_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_1__1__16_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_1__1__16_cbx_1__0__chanx_left_out;
wire [0:64] tile_1__1__16_cby_1__1__chany_top_out;
wire [0:0] tile_1__1__16_ccff_tail;
wire [0:0] tile_1__1__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__1__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__1__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__1__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__1__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__1__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__1__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__1__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__1__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__1__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__1__16_sb_1__0__chanx_right_out;
wire [0:0] tile_1__1__1_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_1__1__1_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_1__1__1_cbx_1__0__chanx_left_out;
wire [0:64] tile_1__1__1_cby_1__1__chany_top_out;
wire [0:0] tile_1__1__1_ccff_tail;
wire [0:0] tile_1__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__1__1_sb_1__0__chanx_right_out;
wire [0:0] tile_1__1__2_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_1__1__2_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_1__1__2_cbx_1__0__chanx_left_out;
wire [0:64] tile_1__1__2_cby_1__1__chany_top_out;
wire [0:0] tile_1__1__2_ccff_tail;
wire [0:0] tile_1__1__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__1__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__1__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__1__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__1__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__1__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__1__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__1__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__1__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__1__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__1__2_sb_1__0__chanx_right_out;
wire [0:0] tile_1__1__3_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_1__1__3_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_1__1__3_cbx_1__0__chanx_left_out;
wire [0:64] tile_1__1__3_cby_1__1__chany_top_out;
wire [0:0] tile_1__1__3_ccff_tail;
wire [0:0] tile_1__1__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__1__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__1__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__1__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__1__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__1__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__1__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__1__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__1__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__1__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__1__3_sb_1__0__chanx_right_out;
wire [0:0] tile_1__1__4_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_1__1__4_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_1__1__4_cbx_1__0__chanx_left_out;
wire [0:64] tile_1__1__4_cby_1__1__chany_top_out;
wire [0:0] tile_1__1__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__1__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__1__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__1__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__1__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__1__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__1__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__1__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__1__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__1__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__1__4_sb_1__0__chanx_right_out;
wire [0:0] tile_1__1__5_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_1__1__5_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_1__1__5_cbx_1__0__chanx_left_out;
wire [0:64] tile_1__1__5_cby_1__1__chany_top_out;
wire [0:0] tile_1__1__5_ccff_tail;
wire [0:0] tile_1__1__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__1__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__1__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__1__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__1__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__1__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__1__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__1__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__1__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__1__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__1__5_sb_1__0__chanx_right_out;
wire [0:0] tile_1__1__6_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_1__1__6_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_1__1__6_cbx_1__0__chanx_left_out;
wire [0:64] tile_1__1__6_cby_1__1__chany_top_out;
wire [0:0] tile_1__1__6_ccff_tail;
wire [0:0] tile_1__1__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__1__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__1__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__1__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__1__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__1__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__1__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__1__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__1__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__1__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__1__6_sb_1__0__chanx_right_out;
wire [0:0] tile_1__1__7_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_1__1__7_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_1__1__7_cbx_1__0__chanx_left_out;
wire [0:64] tile_1__1__7_cby_1__1__chany_top_out;
wire [0:0] tile_1__1__7_ccff_tail;
wire [0:0] tile_1__1__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__1__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__1__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__1__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__1__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__1__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__1__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__1__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__1__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__1__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__1__7_sb_1__0__chanx_right_out;
wire [0:0] tile_1__1__8_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_1__1__8_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_1__1__8_cbx_1__0__chanx_left_out;
wire [0:64] tile_1__1__8_cby_1__1__chany_top_out;
wire [0:0] tile_1__1__8_ccff_tail;
wire [0:0] tile_1__1__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__1__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__1__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__1__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__1__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__1__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__1__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__1__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__1__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__1__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__1__8_sb_1__0__chanx_right_out;
wire [0:0] tile_1__1__9_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_1__1__9_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_1__1__9_cbx_1__0__chanx_left_out;
wire [0:64] tile_1__1__9_cby_1__1__chany_top_out;
wire [0:0] tile_1__1__9_ccff_tail;
wire [0:0] tile_1__1__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__1__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__1__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__1__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__1__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__1__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__1__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__1__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__1__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__1__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__1__9_sb_1__0__chanx_right_out;
wire [0:0] tile_1__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__0_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__0_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__0_ccff_tail;
wire [0:0] tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__0_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__0_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__100_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__100_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__100_ccff_tail;
wire [0:0] tile_1__2__100_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__100_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__100_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__100_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__100_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__100_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__100_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__100_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__100_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__100_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__100_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__100_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__100_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__101_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__101_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__101_ccff_tail;
wire [0:0] tile_1__2__101_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__101_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__101_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__101_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__101_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__101_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__101_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__101_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__101_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__101_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__101_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__101_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__101_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__102_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__102_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__102_ccff_tail;
wire [0:0] tile_1__2__102_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__102_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__102_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__102_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__102_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__102_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__102_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__102_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__102_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__102_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__102_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__102_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__102_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__103_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__103_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__103_ccff_tail;
wire [0:0] tile_1__2__103_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__103_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__103_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__103_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__103_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__103_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__103_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__103_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__103_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__103_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__103_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__103_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__103_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__104_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__104_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__104_ccff_tail;
wire [0:0] tile_1__2__104_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__104_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__104_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__104_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__104_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__104_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__104_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__104_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__104_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__104_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__104_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__104_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__104_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__105_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__105_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__105_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__105_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__105_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__105_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__105_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__105_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__105_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__105_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__105_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__105_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__105_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__105_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__105_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__106_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__106_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__106_ccff_tail;
wire [0:0] tile_1__2__106_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__106_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__106_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__106_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__106_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__106_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__106_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__106_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__106_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__106_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__106_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__106_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__106_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__107_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__107_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__107_ccff_tail;
wire [0:0] tile_1__2__107_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__107_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__107_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__107_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__107_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__107_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__107_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__107_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__107_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__107_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__107_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__107_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__107_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__108_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__108_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__108_ccff_tail;
wire [0:0] tile_1__2__108_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__108_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__108_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__108_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__108_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__108_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__108_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__108_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__108_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__108_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__108_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__108_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__108_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__109_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__109_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__109_ccff_tail;
wire [0:0] tile_1__2__109_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__109_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__109_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__109_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__109_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__109_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__109_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__109_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__109_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__109_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__109_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__109_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__109_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__10_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__10_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__10_ccff_tail;
wire [0:0] tile_1__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__10_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__10_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__110_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__110_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__110_ccff_tail;
wire [0:0] tile_1__2__110_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__110_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__110_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__110_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__110_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__110_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__110_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__110_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__110_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__110_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__110_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__110_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__110_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__111_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__111_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__111_ccff_tail;
wire [0:0] tile_1__2__111_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__111_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__111_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__111_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__111_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__111_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__111_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__111_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__111_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__111_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__111_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__111_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__111_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__112_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__112_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__112_ccff_tail;
wire [0:0] tile_1__2__112_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__112_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__112_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__112_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__112_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__112_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__112_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__112_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__112_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__112_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__112_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__112_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__112_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__113_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__113_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__113_ccff_tail;
wire [0:0] tile_1__2__113_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__113_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__113_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__113_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__113_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__113_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__113_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__113_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__113_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__113_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__113_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__113_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__113_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__114_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__114_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__114_ccff_tail;
wire [0:0] tile_1__2__114_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__114_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__114_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__114_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__114_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__114_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__114_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__114_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__114_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__114_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__114_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__114_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__114_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__115_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__115_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__115_ccff_tail;
wire [0:0] tile_1__2__115_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__115_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__115_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__115_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__115_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__115_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__115_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__115_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__115_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__115_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__115_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__115_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__115_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__116_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__116_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__116_ccff_tail;
wire [0:0] tile_1__2__116_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__116_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__116_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__116_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__116_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__116_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__116_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__116_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__116_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__116_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__116_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__116_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__116_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__117_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__117_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__117_ccff_tail;
wire [0:0] tile_1__2__117_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__117_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__117_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__117_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__117_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__117_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__117_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__117_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__117_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__117_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__117_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__117_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__117_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__118_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__118_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__118_ccff_tail;
wire [0:0] tile_1__2__118_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__118_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__118_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__118_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__118_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__118_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__118_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__118_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__118_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__118_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__118_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__118_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__118_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__119_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__119_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__119_ccff_tail;
wire [0:0] tile_1__2__119_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__119_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__119_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__119_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__119_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__119_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__119_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__119_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__119_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__119_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__119_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__119_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__119_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__11_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__11_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__11_ccff_tail;
wire [0:0] tile_1__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__11_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__11_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__120_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__120_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__120_ccff_tail;
wire [0:0] tile_1__2__120_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__120_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__120_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__120_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__120_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__120_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__120_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__120_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__120_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__120_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__120_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__120_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__120_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__121_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__121_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__121_ccff_tail;
wire [0:0] tile_1__2__121_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__121_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__121_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__121_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__121_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__121_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__121_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__121_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__121_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__121_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__121_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__121_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__121_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__122_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__122_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__122_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__122_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__122_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__122_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__122_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__122_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__122_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__122_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__122_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__122_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__122_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__122_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__122_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__123_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__123_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__123_ccff_tail;
wire [0:0] tile_1__2__123_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__123_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__123_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__123_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__123_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__123_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__123_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__123_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__123_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__123_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__123_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__123_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__123_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__124_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__124_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__124_ccff_tail;
wire [0:0] tile_1__2__124_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__124_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__124_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__124_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__124_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__124_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__124_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__124_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__124_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__124_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__124_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__124_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__124_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__125_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__125_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__125_ccff_tail;
wire [0:0] tile_1__2__125_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__125_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__125_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__125_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__125_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__125_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__125_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__125_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__125_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__125_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__125_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__125_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__125_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__126_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__126_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__126_ccff_tail;
wire [0:0] tile_1__2__126_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__126_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__126_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__126_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__126_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__126_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__126_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__126_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__126_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__126_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__126_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__126_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__126_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__127_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__127_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__127_ccff_tail;
wire [0:0] tile_1__2__127_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__127_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__127_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__127_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__127_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__127_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__127_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__127_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__127_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__127_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__127_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__127_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__127_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__128_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__128_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__128_ccff_tail;
wire [0:0] tile_1__2__128_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__128_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__128_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__128_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__128_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__128_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__128_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__128_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__128_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__128_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__128_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__128_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__128_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__129_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__129_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__129_ccff_tail;
wire [0:0] tile_1__2__129_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__129_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__129_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__129_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__129_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__129_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__129_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__129_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__129_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__129_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__129_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__129_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__129_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__12_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__12_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__12_ccff_tail;
wire [0:0] tile_1__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__12_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__12_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__130_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__130_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__130_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__130_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__130_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__130_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__130_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__130_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__130_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__130_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__130_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__130_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__130_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__130_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__130_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__131_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__131_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__131_ccff_tail;
wire [0:0] tile_1__2__131_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__131_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__131_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__131_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__131_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__131_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__131_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__131_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__131_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__131_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__131_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__131_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__131_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__132_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__132_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__132_ccff_tail;
wire [0:0] tile_1__2__132_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__132_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__132_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__132_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__132_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__132_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__132_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__132_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__132_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__132_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__132_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__132_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__132_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__133_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__133_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__133_ccff_tail;
wire [0:0] tile_1__2__133_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__133_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__133_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__133_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__133_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__133_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__133_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__133_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__133_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__133_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__133_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__133_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__133_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__134_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__134_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__134_ccff_tail;
wire [0:0] tile_1__2__134_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__134_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__134_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__134_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__134_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__134_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__134_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__134_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__134_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__134_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__134_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__134_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__134_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__135_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__135_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__135_ccff_tail;
wire [0:0] tile_1__2__135_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__135_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__135_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__135_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__135_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__135_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__135_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__135_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__135_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__135_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__135_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__135_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__135_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__136_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__136_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__136_ccff_tail;
wire [0:0] tile_1__2__136_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__136_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__136_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__136_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__136_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__136_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__136_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__136_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__136_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__136_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__136_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__136_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__136_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__137_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__137_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__137_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__137_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__137_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__137_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__137_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__137_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__137_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__137_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__137_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__137_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__137_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__137_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__137_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__138_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__138_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__138_ccff_tail;
wire [0:0] tile_1__2__138_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__138_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__138_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__138_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__138_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__138_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__138_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__138_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__138_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__138_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__138_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__138_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__138_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__139_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__139_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__139_ccff_tail;
wire [0:0] tile_1__2__139_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__139_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__139_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__139_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__139_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__139_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__139_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__139_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__139_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__139_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__139_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__139_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__139_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__13_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__13_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__13_ccff_tail;
wire [0:0] tile_1__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__13_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__13_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__140_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__140_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__140_ccff_tail;
wire [0:0] tile_1__2__140_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__140_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__140_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__140_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__140_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__140_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__140_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__140_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__140_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__140_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__140_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__140_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__140_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__141_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__141_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__141_ccff_tail;
wire [0:0] tile_1__2__141_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__141_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__141_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__141_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__141_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__141_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__141_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__141_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__141_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__141_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__141_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__141_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__141_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__142_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__142_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__142_ccff_tail;
wire [0:0] tile_1__2__142_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__142_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__142_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__142_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__142_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__142_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__142_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__142_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__142_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__142_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__142_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__142_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__142_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__143_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__143_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__143_ccff_tail;
wire [0:0] tile_1__2__143_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__143_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__143_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__143_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__143_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__143_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__143_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__143_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__143_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__143_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__143_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__143_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__143_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__144_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__144_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__144_ccff_tail;
wire [0:0] tile_1__2__144_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__144_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__144_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__144_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__144_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__144_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__144_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__144_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__144_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__144_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__144_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__144_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__144_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__145_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__145_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__145_ccff_tail;
wire [0:0] tile_1__2__145_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__145_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__145_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__145_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__145_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__145_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__145_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__145_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__145_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__145_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__145_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__145_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__145_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__146_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__146_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__146_ccff_tail;
wire [0:0] tile_1__2__146_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__146_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__146_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__146_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__146_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__146_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__146_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__146_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__146_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__146_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__146_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__146_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__146_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__147_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__147_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__147_ccff_tail;
wire [0:0] tile_1__2__147_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__147_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__147_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__147_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__147_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__147_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__147_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__147_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__147_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__147_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__147_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__147_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__147_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__148_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__148_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__148_ccff_tail;
wire [0:0] tile_1__2__148_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__148_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__148_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__148_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__148_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__148_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__148_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__148_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__148_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__148_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__148_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__148_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__148_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__149_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__149_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__149_ccff_tail;
wire [0:0] tile_1__2__149_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__149_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__149_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__149_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__149_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__149_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__149_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__149_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__149_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__149_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__149_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__149_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__149_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__14_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__14_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__14_ccff_tail;
wire [0:0] tile_1__2__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__14_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__14_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__14_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__150_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__150_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__150_ccff_tail;
wire [0:0] tile_1__2__150_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__150_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__150_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__150_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__150_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__150_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__150_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__150_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__150_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__150_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__150_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__150_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__150_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__151_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__151_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__151_ccff_tail;
wire [0:0] tile_1__2__151_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__151_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__151_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__151_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__151_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__151_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__151_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__151_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__151_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__151_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__151_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__151_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__151_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__152_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__152_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__152_ccff_tail;
wire [0:0] tile_1__2__152_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__152_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__152_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__152_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__152_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__152_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__152_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__152_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__152_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__152_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__152_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__152_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__152_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__153_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__153_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__153_ccff_tail;
wire [0:0] tile_1__2__153_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__153_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__153_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__153_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__153_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__153_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__153_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__153_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__153_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__153_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__153_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__153_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__153_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__154_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__154_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__154_ccff_tail;
wire [0:0] tile_1__2__154_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__154_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__154_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__154_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__154_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__154_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__154_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__154_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__154_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__154_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__154_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__154_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__154_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__155_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__155_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__155_ccff_tail;
wire [0:0] tile_1__2__155_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__155_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__155_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__155_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__155_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__155_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__155_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__155_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__155_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__155_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__155_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__155_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__155_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__156_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__156_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__156_ccff_tail;
wire [0:0] tile_1__2__156_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__156_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__156_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__156_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__156_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__156_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__156_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__156_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__156_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__156_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__156_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__156_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__156_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__157_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__157_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__157_ccff_tail;
wire [0:0] tile_1__2__157_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__157_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__157_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__157_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__157_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__157_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__157_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__157_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__157_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__157_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__157_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__157_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__157_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__158_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__158_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__158_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__158_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__158_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__158_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__158_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__158_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__158_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__158_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__158_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__158_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__158_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__158_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__158_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__159_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__159_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__159_ccff_tail;
wire [0:0] tile_1__2__159_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__159_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__159_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__159_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__159_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__159_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__159_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__159_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__159_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__159_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__159_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__159_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__159_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__15_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__15_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__15_ccff_tail;
wire [0:0] tile_1__2__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__15_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__15_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__15_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__160_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__160_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__160_ccff_tail;
wire [0:0] tile_1__2__160_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__160_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__160_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__160_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__160_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__160_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__160_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__160_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__160_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__160_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__160_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__160_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__160_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__161_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__161_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__161_ccff_tail;
wire [0:0] tile_1__2__161_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__161_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__161_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__161_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__161_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__161_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__161_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__161_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__161_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__161_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__161_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__161_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__161_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__162_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__162_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__162_ccff_tail;
wire [0:0] tile_1__2__162_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__162_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__162_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__162_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__162_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__162_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__162_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__162_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__162_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__162_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__162_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__162_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__162_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__163_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__163_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__163_ccff_tail;
wire [0:0] tile_1__2__163_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__163_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__163_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__163_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__163_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__163_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__163_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__163_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__163_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__163_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__163_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__163_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__163_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__164_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__164_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__164_ccff_tail;
wire [0:0] tile_1__2__164_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__164_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__164_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__164_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__164_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__164_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__164_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__164_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__164_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__164_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__164_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__164_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__164_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__165_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__165_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__165_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__165_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__165_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__165_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__165_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__165_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__165_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__165_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__165_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__165_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__165_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__165_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__165_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__166_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__166_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__166_ccff_tail;
wire [0:0] tile_1__2__166_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__166_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__166_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__166_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__166_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__166_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__166_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__166_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__166_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__166_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__166_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__166_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__166_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__167_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__167_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__167_ccff_tail;
wire [0:0] tile_1__2__167_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__167_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__167_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__167_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__167_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__167_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__167_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__167_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__167_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__167_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__167_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__167_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__167_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__168_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__168_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__168_ccff_tail;
wire [0:0] tile_1__2__168_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__168_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__168_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__168_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__168_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__168_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__168_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__168_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__168_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__168_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__168_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__168_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__168_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__169_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__169_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__169_ccff_tail;
wire [0:0] tile_1__2__169_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__169_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__169_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__169_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__169_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__169_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__169_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__169_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__169_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__169_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__169_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__169_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__169_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__16_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__16_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__16_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__16_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__16_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__170_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__170_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__170_ccff_tail;
wire [0:0] tile_1__2__170_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__170_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__170_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__170_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__170_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__170_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__170_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__170_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__170_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__170_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__170_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__170_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__170_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__171_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__171_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__171_ccff_tail;
wire [0:0] tile_1__2__171_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__171_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__171_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__171_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__171_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__171_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__171_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__171_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__171_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__171_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__171_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__171_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__171_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__172_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__172_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__172_ccff_tail;
wire [0:0] tile_1__2__172_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__172_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__172_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__172_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__172_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__172_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__172_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__172_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__172_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__172_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__172_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__172_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__172_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__173_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__173_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__173_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__173_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__173_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__173_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__173_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__173_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__173_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__173_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__173_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__173_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__173_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__173_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__173_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__174_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__174_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__174_ccff_tail;
wire [0:0] tile_1__2__174_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__174_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__174_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__174_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__174_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__174_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__174_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__174_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__174_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__174_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__174_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__174_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__174_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__175_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__175_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__175_ccff_tail;
wire [0:0] tile_1__2__175_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__175_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__175_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__175_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__175_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__175_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__175_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__175_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__175_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__175_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__175_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__175_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__175_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__176_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__176_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__176_ccff_tail;
wire [0:0] tile_1__2__176_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__176_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__176_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__176_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__176_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__176_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__176_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__176_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__176_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__176_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__176_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__176_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__176_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__177_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__177_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__177_ccff_tail;
wire [0:0] tile_1__2__177_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__177_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__177_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__177_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__177_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__177_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__177_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__177_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__177_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__177_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__177_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__177_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__177_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__178_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__178_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__178_ccff_tail;
wire [0:0] tile_1__2__178_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__178_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__178_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__178_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__178_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__178_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__178_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__178_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__178_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__178_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__178_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__178_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__178_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__179_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__179_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__179_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__179_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__179_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__179_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__179_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__179_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__179_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__179_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__179_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__179_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__179_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__179_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__179_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__17_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__17_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__17_ccff_tail;
wire [0:0] tile_1__2__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__17_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__17_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__17_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__180_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__180_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__180_ccff_tail;
wire [0:0] tile_1__2__180_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__180_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__180_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__180_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__180_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__180_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__180_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__180_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__180_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__180_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__180_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__180_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__180_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__181_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__181_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__181_ccff_tail;
wire [0:0] tile_1__2__181_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__181_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__181_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__181_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__181_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__181_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__181_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__181_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__181_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__181_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__181_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__181_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__181_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__182_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__182_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__182_ccff_tail;
wire [0:0] tile_1__2__182_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__182_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__182_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__182_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__182_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__182_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__182_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__182_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__182_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__182_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__182_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__182_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__182_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__183_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__183_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__183_ccff_tail;
wire [0:0] tile_1__2__183_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__183_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__183_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__183_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__183_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__183_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__183_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__183_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__183_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__183_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__183_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__183_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__183_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__184_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__184_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__184_ccff_tail;
wire [0:0] tile_1__2__184_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__184_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__184_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__184_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__184_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__184_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__184_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__184_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__184_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__184_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__184_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__184_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__184_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__185_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__185_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__185_ccff_tail;
wire [0:0] tile_1__2__185_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__185_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__185_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__185_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__185_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__185_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__185_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__185_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__185_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__185_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__185_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__185_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__185_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__186_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__186_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__186_ccff_tail;
wire [0:0] tile_1__2__186_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__186_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__186_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__186_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__186_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__186_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__186_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__186_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__186_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__186_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__186_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__186_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__186_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__18_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__18_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__18_ccff_tail;
wire [0:0] tile_1__2__18_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__18_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__18_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__18_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__18_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__18_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__18_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__18_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__18_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__18_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__18_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__18_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__18_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__19_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__19_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__19_ccff_tail;
wire [0:0] tile_1__2__19_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__19_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__19_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__19_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__19_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__19_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__19_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__19_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__19_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__19_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__19_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__19_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__19_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__1_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__1_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__1_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__1_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__20_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__20_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__20_ccff_tail;
wire [0:0] tile_1__2__20_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__20_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__20_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__20_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__20_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__20_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__20_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__20_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__20_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__20_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__20_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__20_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__20_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__21_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__21_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__21_ccff_tail;
wire [0:0] tile_1__2__21_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__21_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__21_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__21_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__21_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__21_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__21_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__21_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__21_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__21_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__21_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__21_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__21_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__22_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__22_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__22_ccff_tail;
wire [0:0] tile_1__2__22_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__22_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__22_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__22_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__22_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__22_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__22_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__22_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__22_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__22_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__22_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__22_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__22_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__23_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__23_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__23_ccff_tail;
wire [0:0] tile_1__2__23_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__23_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__23_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__23_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__23_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__23_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__23_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__23_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__23_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__23_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__23_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__23_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__23_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__24_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__24_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__24_ccff_tail;
wire [0:0] tile_1__2__24_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__24_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__24_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__24_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__24_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__24_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__24_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__24_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__24_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__24_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__24_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__24_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__24_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__25_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__25_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__25_ccff_tail;
wire [0:0] tile_1__2__25_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__25_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__25_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__25_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__25_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__25_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__25_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__25_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__25_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__25_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__25_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__25_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__25_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__26_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__26_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__26_ccff_tail;
wire [0:0] tile_1__2__26_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__26_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__26_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__26_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__26_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__26_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__26_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__26_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__26_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__26_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__26_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__26_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__26_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__27_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__27_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__27_ccff_tail;
wire [0:0] tile_1__2__27_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__27_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__27_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__27_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__27_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__27_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__27_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__27_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__27_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__27_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__27_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__27_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__27_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__28_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__28_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__28_ccff_tail;
wire [0:0] tile_1__2__28_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__28_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__28_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__28_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__28_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__28_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__28_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__28_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__28_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__28_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__28_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__28_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__28_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__29_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__29_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__29_ccff_tail;
wire [0:0] tile_1__2__29_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__29_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__29_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__29_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__29_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__29_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__29_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__29_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__29_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__29_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__29_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__29_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__29_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__2_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__2_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__2_ccff_tail;
wire [0:0] tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__2_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__2_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__30_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__30_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__30_ccff_tail;
wire [0:0] tile_1__2__30_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__30_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__30_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__30_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__30_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__30_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__30_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__30_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__30_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__30_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__30_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__30_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__30_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__31_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__31_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__31_ccff_tail;
wire [0:0] tile_1__2__31_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__31_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__31_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__31_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__31_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__31_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__31_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__31_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__31_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__31_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__31_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__31_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__31_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__32_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__32_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__32_ccff_tail;
wire [0:0] tile_1__2__32_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__32_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__32_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__32_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__32_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__32_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__32_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__32_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__32_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__32_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__32_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__32_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__32_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__33_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__33_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__33_ccff_tail;
wire [0:0] tile_1__2__33_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__33_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__33_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__33_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__33_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__33_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__33_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__33_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__33_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__33_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__33_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__33_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__33_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__34_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__34_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__34_ccff_tail;
wire [0:0] tile_1__2__34_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__34_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__34_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__34_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__34_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__34_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__34_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__34_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__34_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__34_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__34_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__34_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__34_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__35_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__35_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__35_ccff_tail;
wire [0:0] tile_1__2__35_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__35_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__35_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__35_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__35_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__35_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__35_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__35_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__35_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__35_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__35_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__35_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__35_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__36_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__36_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__36_ccff_tail;
wire [0:0] tile_1__2__36_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__36_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__36_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__36_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__36_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__36_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__36_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__36_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__36_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__36_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__36_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__36_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__36_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__37_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__37_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__37_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__37_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__37_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__37_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__37_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__37_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__37_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__37_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__37_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__37_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__37_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__37_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__37_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__38_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__38_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__38_ccff_tail;
wire [0:0] tile_1__2__38_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__38_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__38_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__38_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__38_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__38_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__38_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__38_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__38_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__38_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__38_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__38_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__38_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__39_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__39_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__39_ccff_tail;
wire [0:0] tile_1__2__39_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__39_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__39_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__39_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__39_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__39_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__39_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__39_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__39_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__39_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__39_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__39_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__39_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__3_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__3_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__3_ccff_tail;
wire [0:0] tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__3_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__3_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__40_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__40_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__40_ccff_tail;
wire [0:0] tile_1__2__40_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__40_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__40_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__40_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__40_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__40_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__40_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__40_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__40_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__40_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__40_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__40_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__40_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__41_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__41_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__41_ccff_tail;
wire [0:0] tile_1__2__41_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__41_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__41_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__41_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__41_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__41_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__41_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__41_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__41_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__41_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__41_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__41_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__41_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__42_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__42_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__42_ccff_tail;
wire [0:0] tile_1__2__42_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__42_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__42_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__42_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__42_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__42_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__42_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__42_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__42_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__42_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__42_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__42_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__42_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__43_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__43_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__43_ccff_tail;
wire [0:0] tile_1__2__43_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__43_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__43_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__43_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__43_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__43_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__43_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__43_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__43_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__43_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__43_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__43_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__43_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__44_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__44_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__44_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__44_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__44_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__44_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__44_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__44_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__44_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__44_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__44_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__44_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__44_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__44_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__44_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__45_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__45_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__45_ccff_tail;
wire [0:0] tile_1__2__45_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__45_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__45_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__45_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__45_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__45_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__45_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__45_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__45_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__45_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__45_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__45_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__45_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__46_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__46_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__46_ccff_tail;
wire [0:0] tile_1__2__46_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__46_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__46_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__46_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__46_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__46_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__46_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__46_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__46_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__46_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__46_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__46_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__46_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__47_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__47_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__47_ccff_tail;
wire [0:0] tile_1__2__47_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__47_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__47_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__47_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__47_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__47_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__47_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__47_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__47_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__47_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__47_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__47_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__47_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__48_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__48_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__48_ccff_tail;
wire [0:0] tile_1__2__48_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__48_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__48_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__48_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__48_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__48_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__48_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__48_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__48_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__48_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__48_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__48_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__48_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__49_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__49_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__49_ccff_tail;
wire [0:0] tile_1__2__49_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__49_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__49_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__49_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__49_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__49_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__49_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__49_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__49_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__49_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__49_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__49_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__49_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__4_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__4_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__4_ccff_tail;
wire [0:0] tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__4_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__4_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__50_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__50_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__50_ccff_tail;
wire [0:0] tile_1__2__50_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__50_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__50_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__50_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__50_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__50_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__50_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__50_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__50_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__50_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__50_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__50_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__50_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__51_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__51_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__51_ccff_tail;
wire [0:0] tile_1__2__51_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__51_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__51_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__51_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__51_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__51_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__51_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__51_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__51_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__51_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__51_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__51_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__51_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__52_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__52_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__52_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__52_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__52_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__52_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__52_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__52_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__52_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__52_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__52_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__52_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__52_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__52_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__52_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__53_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__53_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__53_ccff_tail;
wire [0:0] tile_1__2__53_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__53_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__53_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__53_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__53_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__53_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__53_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__53_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__53_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__53_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__53_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__53_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__53_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__54_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__54_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__54_ccff_tail;
wire [0:0] tile_1__2__54_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__54_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__54_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__54_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__54_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__54_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__54_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__54_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__54_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__54_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__54_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__54_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__54_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__55_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__55_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__55_ccff_tail;
wire [0:0] tile_1__2__55_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__55_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__55_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__55_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__55_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__55_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__55_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__55_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__55_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__55_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__55_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__55_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__55_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__56_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__56_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__56_ccff_tail;
wire [0:0] tile_1__2__56_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__56_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__56_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__56_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__56_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__56_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__56_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__56_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__56_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__56_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__56_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__56_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__56_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__57_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__57_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__57_ccff_tail;
wire [0:0] tile_1__2__57_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__57_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__57_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__57_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__57_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__57_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__57_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__57_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__57_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__57_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__57_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__57_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__57_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__58_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__58_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__58_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__58_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__58_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__58_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__58_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__58_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__58_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__58_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__58_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__58_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__58_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__58_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__58_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__59_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__59_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__59_ccff_tail;
wire [0:0] tile_1__2__59_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__59_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__59_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__59_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__59_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__59_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__59_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__59_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__59_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__59_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__59_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__59_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__59_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__5_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__5_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__5_ccff_tail;
wire [0:0] tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__5_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__5_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__60_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__60_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__60_ccff_tail;
wire [0:0] tile_1__2__60_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__60_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__60_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__60_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__60_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__60_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__60_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__60_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__60_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__60_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__60_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__60_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__60_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__61_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__61_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__61_ccff_tail;
wire [0:0] tile_1__2__61_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__61_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__61_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__61_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__61_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__61_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__61_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__61_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__61_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__61_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__61_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__61_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__61_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__62_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__62_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__62_ccff_tail;
wire [0:0] tile_1__2__62_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__62_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__62_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__62_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__62_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__62_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__62_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__62_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__62_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__62_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__62_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__62_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__62_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__63_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__63_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__63_ccff_tail;
wire [0:0] tile_1__2__63_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__63_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__63_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__63_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__63_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__63_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__63_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__63_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__63_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__63_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__63_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__63_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__63_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__64_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__64_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__64_ccff_tail;
wire [0:0] tile_1__2__64_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__64_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__64_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__64_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__64_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__64_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__64_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__64_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__64_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__64_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__64_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__64_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__64_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__65_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__65_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__65_ccff_tail;
wire [0:0] tile_1__2__65_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__65_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__65_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__65_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__65_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__65_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__65_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__65_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__65_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__65_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__65_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__65_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__65_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__66_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__66_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__66_ccff_tail;
wire [0:0] tile_1__2__66_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__66_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__66_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__66_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__66_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__66_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__66_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__66_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__66_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__66_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__66_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__66_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__66_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__67_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__67_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__67_ccff_tail;
wire [0:0] tile_1__2__67_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__67_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__67_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__67_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__67_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__67_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__67_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__67_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__67_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__67_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__67_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__67_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__67_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__68_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__68_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__68_ccff_tail;
wire [0:0] tile_1__2__68_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__68_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__68_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__68_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__68_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__68_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__68_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__68_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__68_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__68_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__68_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__68_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__68_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__69_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__69_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__69_ccff_tail;
wire [0:0] tile_1__2__69_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__69_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__69_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__69_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__69_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__69_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__69_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__69_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__69_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__69_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__69_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__69_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__69_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__6_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__6_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__6_ccff_tail;
wire [0:0] tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__6_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__6_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__70_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__70_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__70_ccff_tail;
wire [0:0] tile_1__2__70_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__70_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__70_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__70_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__70_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__70_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__70_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__70_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__70_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__70_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__70_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__70_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__70_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__71_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__71_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__71_ccff_tail;
wire [0:0] tile_1__2__71_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__71_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__71_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__71_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__71_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__71_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__71_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__71_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__71_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__71_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__71_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__71_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__71_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__72_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__72_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__72_ccff_tail;
wire [0:0] tile_1__2__72_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__72_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__72_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__72_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__72_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__72_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__72_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__72_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__72_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__72_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__72_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__72_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__72_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__73_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__73_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__73_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__73_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__73_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__73_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__73_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__73_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__73_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__73_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__73_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__73_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__73_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__73_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__73_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__74_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__74_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__74_ccff_tail;
wire [0:0] tile_1__2__74_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__74_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__74_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__74_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__74_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__74_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__74_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__74_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__74_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__74_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__74_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__74_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__74_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__75_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__75_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__75_ccff_tail;
wire [0:0] tile_1__2__75_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__75_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__75_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__75_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__75_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__75_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__75_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__75_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__75_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__75_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__75_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__75_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__75_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__76_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__76_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__76_ccff_tail;
wire [0:0] tile_1__2__76_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__76_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__76_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__76_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__76_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__76_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__76_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__76_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__76_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__76_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__76_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__76_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__76_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__77_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__77_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__77_ccff_tail;
wire [0:0] tile_1__2__77_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__77_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__77_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__77_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__77_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__77_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__77_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__77_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__77_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__77_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__77_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__77_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__77_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__78_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__78_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__78_ccff_tail;
wire [0:0] tile_1__2__78_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__78_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__78_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__78_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__78_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__78_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__78_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__78_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__78_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__78_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__78_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__78_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__78_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__79_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__79_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__79_ccff_tail;
wire [0:0] tile_1__2__79_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__79_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__79_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__79_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__79_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__79_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__79_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__79_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__79_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__79_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__79_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__79_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__79_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__7_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__7_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__7_ccff_tail;
wire [0:0] tile_1__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__7_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__7_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__80_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__80_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__80_ccff_tail;
wire [0:0] tile_1__2__80_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__80_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__80_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__80_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__80_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__80_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__80_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__80_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__80_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__80_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__80_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__80_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__80_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__81_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__81_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__81_ccff_tail;
wire [0:0] tile_1__2__81_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__81_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__81_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__81_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__81_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__81_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__81_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__81_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__81_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__81_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__81_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__81_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__81_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__82_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__82_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__82_ccff_tail;
wire [0:0] tile_1__2__82_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__82_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__82_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__82_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__82_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__82_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__82_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__82_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__82_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__82_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__82_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__82_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__82_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__83_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__83_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__83_ccff_tail;
wire [0:0] tile_1__2__83_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__83_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__83_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__83_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__83_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__83_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__83_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__83_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__83_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__83_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__83_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__83_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__83_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__84_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__84_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__84_ccff_tail;
wire [0:0] tile_1__2__84_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__84_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__84_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__84_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__84_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__84_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__84_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__84_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__84_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__84_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__84_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__84_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__84_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__85_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__85_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__85_ccff_tail;
wire [0:0] tile_1__2__85_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__85_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__85_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__85_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__85_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__85_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__85_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__85_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__85_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__85_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__85_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__85_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__85_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__86_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__86_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__86_ccff_tail;
wire [0:0] tile_1__2__86_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__86_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__86_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__86_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__86_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__86_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__86_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__86_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__86_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__86_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__86_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__86_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__86_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__87_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__87_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__87_ccff_tail;
wire [0:0] tile_1__2__87_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__87_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__87_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__87_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__87_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__87_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__87_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__87_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__87_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__87_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__87_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__87_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__87_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__88_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__88_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__88_ccff_tail;
wire [0:0] tile_1__2__88_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__88_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__88_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__88_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__88_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__88_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__88_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__88_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__88_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__88_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__88_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__88_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__88_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__89_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__89_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__89_ccff_tail;
wire [0:0] tile_1__2__89_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__89_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__89_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__89_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__89_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__89_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__89_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__89_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__89_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__89_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__89_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__89_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__89_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__8_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__8_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__8_ccff_tail;
wire [0:0] tile_1__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__8_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__8_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__90_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__90_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__90_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__90_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__90_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__90_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__90_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__90_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__90_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__90_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__90_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__90_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__90_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__90_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__90_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__91_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__91_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__91_ccff_tail;
wire [0:0] tile_1__2__91_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__91_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__91_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__91_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__91_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__91_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__91_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__91_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__91_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__91_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__91_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__91_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__91_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__92_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__92_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__92_ccff_tail;
wire [0:0] tile_1__2__92_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__92_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__92_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__92_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__92_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__92_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__92_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__92_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__92_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__92_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__92_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__92_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__92_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__93_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__93_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__93_ccff_tail;
wire [0:0] tile_1__2__93_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__93_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__93_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__93_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__93_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__93_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__93_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__93_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__93_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__93_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__93_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__93_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__93_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__94_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__94_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__94_ccff_tail;
wire [0:0] tile_1__2__94_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__94_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__94_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__94_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__94_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__94_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__94_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__94_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__94_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__94_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__94_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__94_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__94_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__95_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__95_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__95_ccff_tail;
wire [0:0] tile_1__2__95_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__95_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__95_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__95_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__95_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__95_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__95_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__95_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__95_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__95_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__95_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__95_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__95_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__96_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__96_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__96_ccff_tail;
wire [0:0] tile_1__2__96_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__96_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__96_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__96_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__96_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__96_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__96_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__96_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__96_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__96_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__96_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__96_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__96_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__97_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__97_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__97_ccff_tail;
wire [0:0] tile_1__2__97_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__97_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__97_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__97_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__97_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__97_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__97_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__97_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__97_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__97_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__97_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__97_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__97_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__98_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__98_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__98_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__98_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__98_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__98_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__98_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__98_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__98_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__98_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__98_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__98_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__98_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__98_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__98_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__99_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__99_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__99_ccff_tail;
wire [0:0] tile_1__2__99_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__99_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__99_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__99_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__99_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__99_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__99_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__99_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__99_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__99_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__99_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__99_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__99_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__9_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__9_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__9_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__9_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__0_cbx_1__4__chanx_left_out;
wire [0:0] tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__0_cby_2__5__chany_top_out;
wire [0:0] tile_1__5__0_ccff_tail;
wire [0:0] tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_1__5__0_sb_1__4__chany_bottom_out;
wire [0:64] tile_1__5__0_sb_2__4__chanx_right_out;
wire [0:64] tile_1__5__0_sb_2__4__chany_bottom_out;
wire [0:0] tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__10_cbx_1__4__chanx_left_out;
wire [0:0] tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__10_cby_2__5__chany_top_out;
wire [0:0] tile_1__5__10_ccff_tail;
wire [0:0] tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_1__5__10_sb_1__4__chany_bottom_out;
wire [0:64] tile_1__5__10_sb_2__4__chanx_right_out;
wire [0:64] tile_1__5__10_sb_2__4__chany_bottom_out;
wire [0:0] tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__11_cbx_1__4__chanx_left_out;
wire [0:0] tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__11_cby_2__5__chany_top_out;
wire [0:0] tile_1__5__11_ccff_tail;
wire [0:0] tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_1__5__11_sb_1__4__chany_bottom_out;
wire [0:64] tile_1__5__11_sb_2__4__chanx_right_out;
wire [0:64] tile_1__5__11_sb_2__4__chany_bottom_out;
wire [0:0] tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__12_cbx_1__4__chanx_left_out;
wire [0:0] tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__12_cby_2__5__chany_top_out;
wire [0:0] tile_1__5__12_ccff_tail;
wire [0:0] tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_1__5__12_sb_1__4__chany_bottom_out;
wire [0:64] tile_1__5__12_sb_2__4__chanx_right_out;
wire [0:64] tile_1__5__12_sb_2__4__chany_bottom_out;
wire [0:0] tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__13_cbx_1__4__chanx_left_out;
wire [0:0] tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__13_cby_2__5__chany_top_out;
wire [0:0] tile_1__5__13_ccff_tail;
wire [0:0] tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_1__5__13_sb_1__4__chany_bottom_out;
wire [0:64] tile_1__5__13_sb_2__4__chanx_right_out;
wire [0:64] tile_1__5__13_sb_2__4__chany_bottom_out;
wire [0:0] tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__14_cbx_1__4__chanx_left_out;
wire [0:0] tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__14_cby_2__5__chany_top_out;
wire [0:0] tile_1__5__14_ccff_tail;
wire [0:0] tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_1__5__14_sb_1__4__chany_bottom_out;
wire [0:64] tile_1__5__14_sb_2__4__chanx_right_out;
wire [0:64] tile_1__5__14_sb_2__4__chany_bottom_out;
wire [0:0] tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__15_cbx_1__4__chanx_left_out;
wire [0:0] tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__15_cby_2__5__chany_top_out;
wire [0:0] tile_1__5__15_ccff_tail;
wire [0:0] tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_1__5__15_sb_1__4__chany_bottom_out;
wire [0:64] tile_1__5__15_sb_2__4__chanx_right_out;
wire [0:64] tile_1__5__15_sb_2__4__chany_bottom_out;
wire [0:0] tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__1_cbx_1__4__chanx_left_out;
wire [0:0] tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__1_cby_2__5__chany_top_out;
wire [0:0] tile_1__5__1_ccff_tail;
wire [0:0] tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_1__5__1_sb_1__4__chany_bottom_out;
wire [0:64] tile_1__5__1_sb_2__4__chanx_right_out;
wire [0:64] tile_1__5__1_sb_2__4__chany_bottom_out;
wire [0:0] tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__2_cbx_1__4__chanx_left_out;
wire [0:0] tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__2_cby_2__5__chany_top_out;
wire [0:0] tile_1__5__2_ccff_tail;
wire [0:0] tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_1__5__2_sb_1__4__chany_bottom_out;
wire [0:64] tile_1__5__2_sb_2__4__chanx_right_out;
wire [0:64] tile_1__5__2_sb_2__4__chany_bottom_out;
wire [0:0] tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__3_cbx_1__4__chanx_left_out;
wire [0:0] tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__3_cby_2__5__chany_top_out;
wire [0:0] tile_1__5__3_ccff_tail;
wire [0:0] tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_1__5__3_sb_1__4__chany_bottom_out;
wire [0:64] tile_1__5__3_sb_2__4__chanx_right_out;
wire [0:64] tile_1__5__3_sb_2__4__chany_bottom_out;
wire [0:0] tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__4_cbx_1__4__chanx_left_out;
wire [0:0] tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__4_cby_2__5__chany_top_out;
wire [0:0] tile_1__5__4_ccff_tail;
wire [0:0] tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_1__5__4_sb_1__4__chany_bottom_out;
wire [0:64] tile_1__5__4_sb_2__4__chanx_right_out;
wire [0:64] tile_1__5__4_sb_2__4__chany_bottom_out;
wire [0:0] tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__5_cbx_1__4__chanx_left_out;
wire [0:0] tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__5_cby_2__5__chany_top_out;
wire [0:0] tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_1__5__5_sb_1__4__chany_bottom_out;
wire [0:64] tile_1__5__5_sb_2__4__chanx_right_out;
wire [0:64] tile_1__5__5_sb_2__4__chany_bottom_out;
wire [0:0] tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__6_cbx_1__4__chanx_left_out;
wire [0:0] tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__6_cby_2__5__chany_top_out;
wire [0:0] tile_1__5__6_ccff_tail;
wire [0:0] tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_1__5__6_sb_1__4__chany_bottom_out;
wire [0:64] tile_1__5__6_sb_2__4__chanx_right_out;
wire [0:64] tile_1__5__6_sb_2__4__chany_bottom_out;
wire [0:0] tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__7_cbx_1__4__chanx_left_out;
wire [0:0] tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__7_cby_2__5__chany_top_out;
wire [0:0] tile_1__5__7_ccff_tail;
wire [0:0] tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_1__5__7_sb_1__4__chany_bottom_out;
wire [0:64] tile_1__5__7_sb_2__4__chanx_right_out;
wire [0:64] tile_1__5__7_sb_2__4__chany_bottom_out;
wire [0:0] tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__8_cbx_1__4__chanx_left_out;
wire [0:0] tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__8_cby_2__5__chany_top_out;
wire [0:0] tile_1__5__8_ccff_tail;
wire [0:0] tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_1__5__8_sb_1__4__chany_bottom_out;
wire [0:64] tile_1__5__8_sb_2__4__chanx_right_out;
wire [0:64] tile_1__5__8_sb_2__4__chany_bottom_out;
wire [0:0] tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__9_cbx_1__4__chanx_left_out;
wire [0:0] tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__5__9_cby_2__5__chany_top_out;
wire [0:0] tile_1__5__9_ccff_tail;
wire [0:0] tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_1__5__9_sb_1__4__chany_bottom_out;
wire [0:64] tile_1__5__9_sb_2__4__chanx_right_out;
wire [0:64] tile_1__5__9_sb_2__4__chany_bottom_out;
wire [0:0] tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_1__6__0_cbx_1__5__chanx_left_out;
wire [0:64] tile_1__6__0_cby_1__6__chany_top_out;
wire [0:0] tile_1__6__0_ccff_tail;
wire [0:0] tile_1__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__6__0_sb_1__5__chanx_right_out;
wire [0:0] tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_1__6__10_cbx_1__5__chanx_left_out;
wire [0:64] tile_1__6__10_cby_1__6__chany_top_out;
wire [0:0] tile_1__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__6__10_sb_1__5__chanx_right_out;
wire [0:0] tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_1__6__11_cbx_1__5__chanx_left_out;
wire [0:64] tile_1__6__11_cby_1__6__chany_top_out;
wire [0:0] tile_1__6__11_ccff_tail;
wire [0:0] tile_1__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__6__11_sb_1__5__chanx_right_out;
wire [0:0] tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_1__6__12_cbx_1__5__chanx_left_out;
wire [0:64] tile_1__6__12_cby_1__6__chany_top_out;
wire [0:0] tile_1__6__12_ccff_tail;
wire [0:0] tile_1__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__6__12_sb_1__5__chanx_right_out;
wire [0:0] tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_1__6__13_cbx_1__5__chanx_left_out;
wire [0:64] tile_1__6__13_cby_1__6__chany_top_out;
wire [0:0] tile_1__6__13_ccff_tail;
wire [0:0] tile_1__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__6__13_sb_1__5__chanx_right_out;
wire [0:0] tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_1__6__14_cbx_1__5__chanx_left_out;
wire [0:64] tile_1__6__14_cby_1__6__chany_top_out;
wire [0:0] tile_1__6__14_ccff_tail;
wire [0:0] tile_1__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__6__14_sb_1__5__chanx_right_out;
wire [0:0] tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_1__6__15_cbx_1__5__chanx_left_out;
wire [0:64] tile_1__6__15_cby_1__6__chany_top_out;
wire [0:0] tile_1__6__15_ccff_tail;
wire [0:0] tile_1__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__6__15_sb_1__5__chanx_right_out;
wire [0:0] tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_1__6__16_cbx_1__5__chanx_left_out;
wire [0:64] tile_1__6__16_cby_1__6__chany_top_out;
wire [0:0] tile_1__6__16_ccff_tail;
wire [0:0] tile_1__6__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__6__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__6__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__6__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__6__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__6__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__6__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__6__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__6__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__6__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__6__16_sb_1__5__chanx_right_out;
wire [0:0] tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_1__6__17_cbx_1__5__chanx_left_out;
wire [0:64] tile_1__6__17_cby_1__6__chany_top_out;
wire [0:0] tile_1__6__17_ccff_tail;
wire [0:0] tile_1__6__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__6__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__6__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__6__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__6__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__6__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__6__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__6__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__6__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__6__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__6__17_sb_1__5__chanx_right_out;
wire [0:0] tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_1__6__1_cbx_1__5__chanx_left_out;
wire [0:64] tile_1__6__1_cby_1__6__chany_top_out;
wire [0:0] tile_1__6__1_ccff_tail;
wire [0:0] tile_1__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__6__1_sb_1__5__chanx_right_out;
wire [0:0] tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_1__6__2_cbx_1__5__chanx_left_out;
wire [0:64] tile_1__6__2_cby_1__6__chany_top_out;
wire [0:0] tile_1__6__2_ccff_tail;
wire [0:0] tile_1__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__6__2_sb_1__5__chanx_right_out;
wire [0:0] tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_1__6__3_cbx_1__5__chanx_left_out;
wire [0:64] tile_1__6__3_cby_1__6__chany_top_out;
wire [0:0] tile_1__6__3_ccff_tail;
wire [0:0] tile_1__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__6__3_sb_1__5__chanx_right_out;
wire [0:0] tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_1__6__4_cbx_1__5__chanx_left_out;
wire [0:64] tile_1__6__4_cby_1__6__chany_top_out;
wire [0:0] tile_1__6__4_ccff_tail;
wire [0:0] tile_1__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__6__4_sb_1__5__chanx_right_out;
wire [0:0] tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_1__6__5_cbx_1__5__chanx_left_out;
wire [0:64] tile_1__6__5_cby_1__6__chany_top_out;
wire [0:0] tile_1__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__6__5_sb_1__5__chanx_right_out;
wire [0:0] tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_1__6__6_cbx_1__5__chanx_left_out;
wire [0:64] tile_1__6__6_cby_1__6__chany_top_out;
wire [0:0] tile_1__6__6_ccff_tail;
wire [0:0] tile_1__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__6__6_sb_1__5__chanx_right_out;
wire [0:0] tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_1__6__7_cbx_1__5__chanx_left_out;
wire [0:64] tile_1__6__7_cby_1__6__chany_top_out;
wire [0:0] tile_1__6__7_ccff_tail;
wire [0:0] tile_1__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__6__7_sb_1__5__chanx_right_out;
wire [0:0] tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_1__6__8_cbx_1__5__chanx_left_out;
wire [0:64] tile_1__6__8_cby_1__6__chany_top_out;
wire [0:0] tile_1__6__8_ccff_tail;
wire [0:0] tile_1__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__6__8_sb_1__5__chanx_right_out;
wire [0:0] tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_1__6__9_cbx_1__5__chanx_left_out;
wire [0:64] tile_1__6__9_cby_1__6__chany_top_out;
wire [0:0] tile_1__6__9_ccff_tail;
wire [0:0] tile_1__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__6__9_sb_1__5__chanx_right_out;
wire [0:0] tile_1__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:64] tile_2__11__0_cbx_2__10__chanx_left_out;
wire [0:64] tile_2__11__0_cby_2__11__chany_top_out;
wire [0:0] tile_2__11__0_ccff_tail;
wire [0:0] tile_2__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__11__0_sb_2__10__chanx_right_out;
wire [0:64] tile_2__11__0_sb_2__10__chany_bottom_out;
wire [0:64] tile_2__11__1_cbx_2__10__chanx_left_out;
wire [0:64] tile_2__11__1_cby_2__11__chany_top_out;
wire [0:0] tile_2__11__1_ccff_tail;
wire [0:0] tile_2__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__11__1_sb_2__10__chanx_right_out;
wire [0:64] tile_2__11__1_sb_2__10__chany_bottom_out;
wire [0:64] tile_2__11__2_cbx_2__10__chanx_left_out;
wire [0:64] tile_2__11__2_cby_2__11__chany_top_out;
wire [0:0] tile_2__11__2_ccff_tail;
wire [0:0] tile_2__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__11__2_sb_2__10__chanx_right_out;
wire [0:64] tile_2__11__2_sb_2__10__chany_bottom_out;
wire [0:64] tile_2__11__3_cbx_2__10__chanx_left_out;
wire [0:64] tile_2__11__3_cby_2__11__chany_top_out;
wire [0:0] tile_2__11__3_ccff_tail;
wire [0:0] tile_2__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__11__3_sb_2__10__chanx_right_out;
wire [0:64] tile_2__11__3_sb_2__10__chany_bottom_out;
wire [0:64] tile_2__11__4_cbx_2__10__chanx_left_out;
wire [0:64] tile_2__11__4_cby_2__11__chany_top_out;
wire [0:0] tile_2__11__4_ccff_tail;
wire [0:0] tile_2__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__11__4_sb_2__10__chanx_right_out;
wire [0:64] tile_2__11__4_sb_2__10__chany_bottom_out;
wire [0:64] tile_2__11__5_cbx_2__10__chanx_left_out;
wire [0:64] tile_2__11__5_cby_2__11__chany_top_out;
wire [0:0] tile_2__11__5_ccff_tail;
wire [0:0] tile_2__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__11__5_sb_2__10__chanx_right_out;
wire [0:64] tile_2__11__5_sb_2__10__chany_bottom_out;
wire [0:64] tile_2__11__6_cbx_2__10__chanx_left_out;
wire [0:64] tile_2__11__6_cby_2__11__chany_top_out;
wire [0:0] tile_2__11__6_ccff_tail;
wire [0:0] tile_2__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__11__6_sb_2__10__chanx_right_out;
wire [0:64] tile_2__11__6_sb_2__10__chany_bottom_out;
wire [0:64] tile_2__11__7_cbx_2__10__chanx_left_out;
wire [0:64] tile_2__11__7_cby_2__11__chany_top_out;
wire [0:0] tile_2__11__7_ccff_tail;
wire [0:0] tile_2__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__11__7_sb_2__10__chanx_right_out;
wire [0:64] tile_2__11__7_sb_2__10__chany_bottom_out;
wire [0:0] tile_2__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_2__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_2__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_2__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_2__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_2__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:64] tile_2__6__0_cbx_2__5__chanx_left_out;
wire [0:64] tile_2__6__0_cby_2__6__chany_top_out;
wire [0:0] tile_2__6__0_ccff_tail;
wire [0:0] tile_2__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__6__0_sb_2__5__chanx_right_out;
wire [0:64] tile_2__6__0_sb_2__5__chany_bottom_out;
wire [0:64] tile_2__6__10_cbx_2__5__chanx_left_out;
wire [0:64] tile_2__6__10_cby_2__6__chany_top_out;
wire [0:0] tile_2__6__10_ccff_tail;
wire [0:0] tile_2__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__6__10_sb_2__5__chanx_right_out;
wire [0:64] tile_2__6__10_sb_2__5__chany_bottom_out;
wire [0:64] tile_2__6__11_cbx_2__5__chanx_left_out;
wire [0:64] tile_2__6__11_cby_2__6__chany_top_out;
wire [0:0] tile_2__6__11_ccff_tail;
wire [0:0] tile_2__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__6__11_sb_2__5__chanx_right_out;
wire [0:64] tile_2__6__11_sb_2__5__chany_bottom_out;
wire [0:64] tile_2__6__12_cbx_2__5__chanx_left_out;
wire [0:64] tile_2__6__12_cby_2__6__chany_top_out;
wire [0:0] tile_2__6__12_ccff_tail;
wire [0:0] tile_2__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__6__12_sb_2__5__chanx_right_out;
wire [0:64] tile_2__6__12_sb_2__5__chany_bottom_out;
wire [0:64] tile_2__6__13_cbx_2__5__chanx_left_out;
wire [0:64] tile_2__6__13_cby_2__6__chany_top_out;
wire [0:0] tile_2__6__13_ccff_tail;
wire [0:0] tile_2__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__6__13_sb_2__5__chanx_right_out;
wire [0:64] tile_2__6__13_sb_2__5__chany_bottom_out;
wire [0:64] tile_2__6__14_cbx_2__5__chanx_left_out;
wire [0:64] tile_2__6__14_cby_2__6__chany_top_out;
wire [0:0] tile_2__6__14_ccff_tail;
wire [0:0] tile_2__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__6__14_sb_2__5__chanx_right_out;
wire [0:64] tile_2__6__14_sb_2__5__chany_bottom_out;
wire [0:64] tile_2__6__15_cbx_2__5__chanx_left_out;
wire [0:64] tile_2__6__15_cby_2__6__chany_top_out;
wire [0:0] tile_2__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__6__15_sb_2__5__chanx_right_out;
wire [0:64] tile_2__6__15_sb_2__5__chany_bottom_out;
wire [0:64] tile_2__6__1_cbx_2__5__chanx_left_out;
wire [0:64] tile_2__6__1_cby_2__6__chany_top_out;
wire [0:0] tile_2__6__1_ccff_tail;
wire [0:0] tile_2__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__6__1_sb_2__5__chanx_right_out;
wire [0:64] tile_2__6__1_sb_2__5__chany_bottom_out;
wire [0:64] tile_2__6__2_cbx_2__5__chanx_left_out;
wire [0:64] tile_2__6__2_cby_2__6__chany_top_out;
wire [0:0] tile_2__6__2_ccff_tail;
wire [0:0] tile_2__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__6__2_sb_2__5__chanx_right_out;
wire [0:64] tile_2__6__2_sb_2__5__chany_bottom_out;
wire [0:64] tile_2__6__3_cbx_2__5__chanx_left_out;
wire [0:64] tile_2__6__3_cby_2__6__chany_top_out;
wire [0:0] tile_2__6__3_ccff_tail;
wire [0:0] tile_2__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__6__3_sb_2__5__chanx_right_out;
wire [0:64] tile_2__6__3_sb_2__5__chany_bottom_out;
wire [0:64] tile_2__6__4_cbx_2__5__chanx_left_out;
wire [0:64] tile_2__6__4_cby_2__6__chany_top_out;
wire [0:0] tile_2__6__4_ccff_tail;
wire [0:0] tile_2__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__6__4_sb_2__5__chanx_right_out;
wire [0:64] tile_2__6__4_sb_2__5__chany_bottom_out;
wire [0:64] tile_2__6__5_cbx_2__5__chanx_left_out;
wire [0:64] tile_2__6__5_cby_2__6__chany_top_out;
wire [0:0] tile_2__6__5_ccff_tail;
wire [0:0] tile_2__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__6__5_sb_2__5__chanx_right_out;
wire [0:64] tile_2__6__5_sb_2__5__chany_bottom_out;
wire [0:64] tile_2__6__6_cbx_2__5__chanx_left_out;
wire [0:64] tile_2__6__6_cby_2__6__chany_top_out;
wire [0:0] tile_2__6__6_ccff_tail;
wire [0:0] tile_2__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__6__6_sb_2__5__chanx_right_out;
wire [0:64] tile_2__6__6_sb_2__5__chany_bottom_out;
wire [0:64] tile_2__6__7_cbx_2__5__chanx_left_out;
wire [0:64] tile_2__6__7_cby_2__6__chany_top_out;
wire [0:0] tile_2__6__7_ccff_tail;
wire [0:0] tile_2__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__6__7_sb_2__5__chanx_right_out;
wire [0:64] tile_2__6__7_sb_2__5__chany_bottom_out;
wire [0:64] tile_2__6__8_cbx_2__5__chanx_left_out;
wire [0:64] tile_2__6__8_cby_2__6__chany_top_out;
wire [0:0] tile_2__6__8_ccff_tail;
wire [0:0] tile_2__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__6__8_sb_2__5__chanx_right_out;
wire [0:64] tile_2__6__8_sb_2__5__chany_bottom_out;
wire [0:64] tile_2__6__9_cbx_2__5__chanx_left_out;
wire [0:64] tile_2__6__9_cby_2__6__chany_top_out;
wire [0:0] tile_2__6__9_ccff_tail;
wire [0:0] tile_2__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_2__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_2__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_2__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_2__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_2__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_2__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_2__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_2__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_2__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_2__6__9_sb_2__5__chanx_right_out;
wire [0:64] tile_2__6__9_sb_2__5__chany_bottom_out;
wire [0:0] tile_2__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_2__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_3__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_3__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_3__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_3__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_3__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_3__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_3__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_3__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_4__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_4__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_4__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_4__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_4__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_4__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_4__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_4__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_5__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_5__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_5__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_5__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_5__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_5__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_5__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_5__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_6__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_6__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_6__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_6__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_6__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_6__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_6__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_6__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_7__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_7__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_7__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_7__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_7__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_7__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_7__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_7__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_8__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_8__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_8__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_8__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_8__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_8__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_8__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_8__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_9__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_9__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_9__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_9__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_9__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_9__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_9__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_9__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	tile_0__19_ tile_0__19_ (
		.prog_clk(prog_clk),
		.sb_0__18__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__18__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__10_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__18__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__10_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__18__chanx_right_in(tile_1__19__0_cbx_1__18__chanx_left_out[0:64]),
		.sb_0__18__chany_bottom_in(tile_0__2__10_cby_0__2__chany_top_out[0:64]),
		.ccff_head(tile_1__19__0_ccff_tail),
		.sb_0__18__chanx_right_out(tile_0__19__0_sb_0__18__chanx_right_out[0:64]),
		.sb_0__18__chany_bottom_out(tile_0__19__0_sb_0__18__chany_bottom_out[0:64]),
		.ccff_tail(ccff_tail[31]));

	tile_1__19_ tile_1__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[0:1]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[0:1]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[0:1]),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__1_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__1_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__chanx_right_in(tile_1__19__1_cbx_1__18__chanx_left_out[0:64]),
		.sb_1__18__chany_bottom_in(tile_1__2__10_cby_1__2__chany_top_out[0:64]),
		.cbx_1__18__chanx_left_in(tile_0__19__0_sb_0__18__chanx_right_out[0:64]),
		.ccff_head(tile_1__19__1_ccff_tail),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__18__chanx_right_out(tile_1__19__0_sb_1__18__chanx_right_out[0:64]),
		.sb_1__18__chany_bottom_out(tile_1__19__0_sb_1__18__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_1__18__chanx_left_out(tile_1__19__0_cbx_1__18__chanx_left_out[0:64]),
		.ccff_tail(tile_1__19__0_ccff_tail));

	tile_1__19_ tile_2__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[2:3]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[2:3]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[2:3]),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__2_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__2_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__21_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__21_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__21_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__21_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__chanx_right_in(tile_1__19__2_cbx_1__18__chanx_left_out[0:64]),
		.sb_1__18__chany_bottom_in(tile_1__2__21_cby_1__2__chany_top_out[0:64]),
		.cbx_1__18__chanx_left_in(tile_1__19__0_sb_1__18__chanx_right_out[0:64]),
		.ccff_head(tile_1__19__2_ccff_tail),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__18__chanx_right_out(tile_1__19__1_sb_1__18__chanx_right_out[0:64]),
		.sb_1__18__chany_bottom_out(tile_1__19__1_sb_1__18__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__1_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__1_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_1__18__chanx_left_out(tile_1__19__1_cbx_1__18__chanx_left_out[0:64]),
		.ccff_tail(tile_1__19__1_ccff_tail));

	tile_1__19_ tile_3__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[4:5]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[4:5]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[4:5]),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__3_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__3_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__32_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__32_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__32_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__32_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__chanx_right_in(tile_1__19__3_cbx_1__18__chanx_left_out[0:64]),
		.sb_1__18__chany_bottom_in(tile_1__2__32_cby_1__2__chany_top_out[0:64]),
		.cbx_1__18__chanx_left_in(tile_1__19__1_sb_1__18__chanx_right_out[0:64]),
		.ccff_head(tile_1__19__3_ccff_tail),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__18__chanx_right_out(tile_1__19__2_sb_1__18__chanx_right_out[0:64]),
		.sb_1__18__chany_bottom_out(tile_1__19__2_sb_1__18__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__2_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__2_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_1__18__chanx_left_out(tile_1__19__2_cbx_1__18__chanx_left_out[0:64]),
		.ccff_tail(tile_1__19__2_ccff_tail));

	tile_1__19_ tile_4__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[6:7]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[6:7]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[6:7]),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__4_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__4_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__43_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__43_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__43_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__43_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__chanx_right_in(tile_1__19__4_cbx_1__18__chanx_left_out[0:64]),
		.sb_1__18__chany_bottom_in(tile_1__2__43_cby_1__2__chany_top_out[0:64]),
		.cbx_1__18__chanx_left_in(tile_1__19__2_sb_1__18__chanx_right_out[0:64]),
		.ccff_head(tile_1__19__4_ccff_tail),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__18__chanx_right_out(tile_1__19__3_sb_1__18__chanx_right_out[0:64]),
		.sb_1__18__chany_bottom_out(tile_1__19__3_sb_1__18__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__3_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__3_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_1__18__chanx_left_out(tile_1__19__3_cbx_1__18__chanx_left_out[0:64]),
		.ccff_tail(tile_1__19__3_ccff_tail));

	tile_1__19_ tile_5__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[8:9]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[8:9]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[8:9]),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__5_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__5_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__54_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__54_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__54_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__54_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__chanx_right_in(tile_1__19__5_cbx_1__18__chanx_left_out[0:64]),
		.sb_1__18__chany_bottom_in(tile_1__2__54_cby_1__2__chany_top_out[0:64]),
		.cbx_1__18__chanx_left_in(tile_1__19__3_sb_1__18__chanx_right_out[0:64]),
		.ccff_head(tile_1__19__5_ccff_tail),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__18__chanx_right_out(tile_1__19__4_sb_1__18__chanx_right_out[0:64]),
		.sb_1__18__chany_bottom_out(tile_1__19__4_sb_1__18__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__4_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__4_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_1__18__chanx_left_out(tile_1__19__4_cbx_1__18__chanx_left_out[0:64]),
		.ccff_tail(tile_1__19__4_ccff_tail));

	tile_1__19_ tile_6__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[10:11]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[10:11]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[10:11]),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__6_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__6_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__65_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__65_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__65_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__65_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__chanx_right_in(tile_1__19__6_cbx_1__18__chanx_left_out[0:64]),
		.sb_1__18__chany_bottom_in(tile_1__2__65_cby_1__2__chany_top_out[0:64]),
		.cbx_1__18__chanx_left_in(tile_1__19__4_sb_1__18__chanx_right_out[0:64]),
		.ccff_head(tile_1__19__6_ccff_tail),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__18__chanx_right_out(tile_1__19__5_sb_1__18__chanx_right_out[0:64]),
		.sb_1__18__chany_bottom_out(tile_1__19__5_sb_1__18__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__5_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__5_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_1__18__chanx_left_out(tile_1__19__5_cbx_1__18__chanx_left_out[0:64]),
		.ccff_tail(tile_1__19__5_ccff_tail));

	tile_1__19_ tile_7__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[12:13]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[12:13]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[12:13]),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__7_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__7_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__76_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__76_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__76_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__76_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__chanx_right_in(tile_1__19__7_cbx_1__18__chanx_left_out[0:64]),
		.sb_1__18__chany_bottom_in(tile_1__2__76_cby_1__2__chany_top_out[0:64]),
		.cbx_1__18__chanx_left_in(tile_1__19__5_sb_1__18__chanx_right_out[0:64]),
		.ccff_head(tile_1__19__7_ccff_tail),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__18__chanx_right_out(tile_1__19__6_sb_1__18__chanx_right_out[0:64]),
		.sb_1__18__chany_bottom_out(tile_1__19__6_sb_1__18__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__6_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__6_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_1__18__chanx_left_out(tile_1__19__6_cbx_1__18__chanx_left_out[0:64]),
		.ccff_tail(tile_1__19__6_ccff_tail));

	tile_1__19_ tile_8__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[14:15]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[14:15]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[14:15]),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__8_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__8_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__87_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__87_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__87_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__87_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__chanx_right_in(tile_1__19__8_cbx_1__18__chanx_left_out[0:64]),
		.sb_1__18__chany_bottom_in(tile_1__2__87_cby_1__2__chany_top_out[0:64]),
		.cbx_1__18__chanx_left_in(tile_1__19__6_sb_1__18__chanx_right_out[0:64]),
		.ccff_head(tile_1__19__8_ccff_tail),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__18__chanx_right_out(tile_1__19__7_sb_1__18__chanx_right_out[0:64]),
		.sb_1__18__chany_bottom_out(tile_1__19__7_sb_1__18__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__7_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__7_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_1__18__chanx_left_out(tile_1__19__7_cbx_1__18__chanx_left_out[0:64]),
		.ccff_tail(tile_1__19__7_ccff_tail));

	tile_1__19_ tile_9__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[16:17]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[16:17]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[16:17]),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__9_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__9_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__98_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__98_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__98_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__98_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__chanx_right_in(tile_1__19__9_cbx_1__18__chanx_left_out[0:64]),
		.sb_1__18__chany_bottom_in(tile_1__2__98_cby_1__2__chany_top_out[0:64]),
		.cbx_1__18__chanx_left_in(tile_1__19__7_sb_1__18__chanx_right_out[0:64]),
		.ccff_head(tile_1__19__9_ccff_tail),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__18__chanx_right_out(tile_1__19__8_sb_1__18__chanx_right_out[0:64]),
		.sb_1__18__chany_bottom_out(tile_1__19__8_sb_1__18__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__8_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__8_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_1__18__chanx_left_out(tile_1__19__8_cbx_1__18__chanx_left_out[0:64]),
		.ccff_tail(tile_1__19__8_ccff_tail));

	tile_1__19_ tile_10__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[18:19]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[18:19]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[18:19]),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__10_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__10_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__109_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__109_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__109_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__109_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__chanx_right_in(tile_1__19__10_cbx_1__18__chanx_left_out[0:64]),
		.sb_1__18__chany_bottom_in(tile_1__2__109_cby_1__2__chany_top_out[0:64]),
		.cbx_1__18__chanx_left_in(tile_1__19__8_sb_1__18__chanx_right_out[0:64]),
		.ccff_head(tile_1__19__10_ccff_tail),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__18__chanx_right_out(tile_1__19__9_sb_1__18__chanx_right_out[0:64]),
		.sb_1__18__chany_bottom_out(tile_1__19__9_sb_1__18__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__9_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__9_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_1__18__chanx_left_out(tile_1__19__9_cbx_1__18__chanx_left_out[0:64]),
		.ccff_tail(tile_1__19__9_ccff_tail));

	tile_1__19_ tile_11__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[20:21]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[20:21]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[20:21]),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__11_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__11_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__120_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__120_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__120_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__120_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__chanx_right_in(tile_1__19__11_cbx_1__18__chanx_left_out[0:64]),
		.sb_1__18__chany_bottom_in(tile_1__2__120_cby_1__2__chany_top_out[0:64]),
		.cbx_1__18__chanx_left_in(tile_1__19__9_sb_1__18__chanx_right_out[0:64]),
		.ccff_head(tile_1__19__11_ccff_tail),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__18__chanx_right_out(tile_1__19__10_sb_1__18__chanx_right_out[0:64]),
		.sb_1__18__chany_bottom_out(tile_1__19__10_sb_1__18__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__10_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__10_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_1__18__chanx_left_out(tile_1__19__10_cbx_1__18__chanx_left_out[0:64]),
		.ccff_tail(tile_1__19__10_ccff_tail));

	tile_1__19_ tile_12__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[22:23]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[22:23]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[22:23]),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__12_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__12_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__131_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__131_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__131_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__131_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__chanx_right_in(tile_1__19__12_cbx_1__18__chanx_left_out[0:64]),
		.sb_1__18__chany_bottom_in(tile_1__2__131_cby_1__2__chany_top_out[0:64]),
		.cbx_1__18__chanx_left_in(tile_1__19__10_sb_1__18__chanx_right_out[0:64]),
		.ccff_head(tile_1__19__12_ccff_tail),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__18__chanx_right_out(tile_1__19__11_sb_1__18__chanx_right_out[0:64]),
		.sb_1__18__chany_bottom_out(tile_1__19__11_sb_1__18__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__11_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__11_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_1__18__chanx_left_out(tile_1__19__11_cbx_1__18__chanx_left_out[0:64]),
		.ccff_tail(tile_1__19__11_ccff_tail));

	tile_1__19_ tile_13__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[24:25]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[24:25]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[24:25]),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__13_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__13_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__142_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__142_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__142_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__142_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__chanx_right_in(tile_1__19__13_cbx_1__18__chanx_left_out[0:64]),
		.sb_1__18__chany_bottom_in(tile_1__2__142_cby_1__2__chany_top_out[0:64]),
		.cbx_1__18__chanx_left_in(tile_1__19__11_sb_1__18__chanx_right_out[0:64]),
		.ccff_head(tile_1__19__13_ccff_tail),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__18__chanx_right_out(tile_1__19__12_sb_1__18__chanx_right_out[0:64]),
		.sb_1__18__chany_bottom_out(tile_1__19__12_sb_1__18__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__12_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__12_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_1__18__chanx_left_out(tile_1__19__12_cbx_1__18__chanx_left_out[0:64]),
		.ccff_tail(tile_1__19__12_ccff_tail));

	tile_1__19_ tile_14__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[26:27]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[26:27]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[26:27]),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__14_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__14_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__153_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__153_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__153_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__153_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__chanx_right_in(tile_1__19__14_cbx_1__18__chanx_left_out[0:64]),
		.sb_1__18__chany_bottom_in(tile_1__2__153_cby_1__2__chany_top_out[0:64]),
		.cbx_1__18__chanx_left_in(tile_1__19__12_sb_1__18__chanx_right_out[0:64]),
		.ccff_head(tile_1__19__14_ccff_tail),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__18__chanx_right_out(tile_1__19__13_sb_1__18__chanx_right_out[0:64]),
		.sb_1__18__chany_bottom_out(tile_1__19__13_sb_1__18__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__13_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__13_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_1__18__chanx_left_out(tile_1__19__13_cbx_1__18__chanx_left_out[0:64]),
		.ccff_tail(tile_1__19__13_ccff_tail));

	tile_1__19_ tile_15__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[28:29]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[28:29]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[28:29]),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__15_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__15_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__164_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__164_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__164_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__164_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__chanx_right_in(tile_1__19__15_cbx_1__18__chanx_left_out[0:64]),
		.sb_1__18__chany_bottom_in(tile_1__2__164_cby_1__2__chany_top_out[0:64]),
		.cbx_1__18__chanx_left_in(tile_1__19__13_sb_1__18__chanx_right_out[0:64]),
		.ccff_head(tile_1__19__15_ccff_tail),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__18__chanx_right_out(tile_1__19__14_sb_1__18__chanx_right_out[0:64]),
		.sb_1__18__chany_bottom_out(tile_1__19__14_sb_1__18__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__14_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__14_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_1__18__chanx_left_out(tile_1__19__14_cbx_1__18__chanx_left_out[0:64]),
		.ccff_tail(tile_1__19__14_ccff_tail));

	tile_1__19_ tile_16__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[30:31]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[30:31]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[30:31]),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__16_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__16_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__175_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__175_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__175_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__175_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__chanx_right_in(tile_1__19__16_cbx_1__18__chanx_left_out[0:64]),
		.sb_1__18__chany_bottom_in(tile_1__2__175_cby_1__2__chany_top_out[0:64]),
		.cbx_1__18__chanx_left_in(tile_1__19__14_sb_1__18__chanx_right_out[0:64]),
		.ccff_head(tile_1__19__16_ccff_tail),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__18__chanx_right_out(tile_1__19__15_sb_1__18__chanx_right_out[0:64]),
		.sb_1__18__chany_bottom_out(tile_1__19__15_sb_1__18__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__15_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__15_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_1__18__chanx_left_out(tile_1__19__15_cbx_1__18__chanx_left_out[0:64]),
		.ccff_tail(tile_1__19__15_ccff_tail));

	tile_1__19_ tile_17__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[32:33]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[32:33]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[32:33]),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_18__19__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__18__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_18__19__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__186_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__186_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__186_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__186_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__18__chanx_right_in(tile_18__19__0_cbx_18__18__chanx_left_out[0:64]),
		.sb_1__18__chany_bottom_in(tile_1__2__186_cby_1__2__chany_top_out[0:64]),
		.cbx_1__18__chanx_left_in(tile_1__19__15_sb_1__18__chanx_right_out[0:64]),
		.ccff_head(tile_18__19__0_ccff_tail),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__18__chanx_right_out(tile_1__19__16_sb_1__18__chanx_right_out[0:64]),
		.sb_1__18__chany_bottom_out(tile_1__19__16_sb_1__18__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__19__16_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__19__16_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_1__18__chanx_left_out(tile_1__19__16_cbx_1__18__chanx_left_out[0:64]),
		.ccff_tail(tile_1__19__16_ccff_tail));

	tile_18__19_ tile_18__19_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[34:35]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[34:35]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[34:35]),
		.sb_18__18__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__0_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__18__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__0_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_18__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_18__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_18__18__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_18__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_18__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_18__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_18__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_18__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_18__18__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_18__18__chany_bottom_in(tile_18__2__10_cby_18__2__chany_top_out[0:64]),
		.cbx_18__18__chanx_left_in(tile_1__19__16_sb_1__18__chanx_right_out[0:64]),
		.ccff_head(tile_19__1__0_ccff_tail),
		.cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_18__18__chany_bottom_out(tile_18__19__0_sb_18__18__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_18__19__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_18__19__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_18__18__chanx_left_out(tile_18__19__0_cbx_18__18__chanx_left_out[0:64]),
		.ccff_tail(tile_18__19__0_ccff_tail));

	tile_19__1_ tile_19__18_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[36:37]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[36:37]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[36:37]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__10_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__10_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_18__2__10_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__0_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__0_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_19__1__0_ccff_tail));

	tile_19__1_ tile_19__17_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[38:39]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[38:39]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[38:39]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__9_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__9_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_19__1__2_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__1_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__1_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_19__1__1_ccff_tail));

	tile_19__1_ tile_19__16_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[40:41]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[40:41]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[40:41]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__8_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__8_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_18__2__8_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__2_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__2_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_19__1__2_ccff_tail));

	tile_19__1_ tile_19__15_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[42:43]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[42:43]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[42:43]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__6__2_cby_18__6__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__6__2_cby_18__6__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_19__1__4_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__3_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__3_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_19__1__3_ccff_tail));

	tile_19__1_ tile_19__14_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[44:45]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[44:45]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[44:45]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_17__5__1_cby_18__5__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_17__5__1_cby_18__5__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_17__5__1_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__4_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__4_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_19__1__4_ccff_tail));

	tile_19__1_ tile_19__13_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[46:47]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[46:47]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[46:47]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__7_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__7_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_19__1__6_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__5_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__5_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_19__1__5_ccff_tail));

	tile_19__1_ tile_19__12_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[48:49]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[48:49]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[48:49]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__6_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__6_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_18__2__6_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__6_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__6_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_19__1__6_ccff_tail));

	tile_19__1_ tile_19__11_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[50:51]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[50:51]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[50:51]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__6__1_cby_18__6__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__6__1_cby_18__6__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_19__1__8_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__7_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__7_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_19__1__7_ccff_tail));

	tile_19__1_ tile_19__10_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[52:53]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[52:53]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[52:53]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_17__10__0_cby_18__10__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_17__10__0_cby_18__10__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_17__10__0_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__8_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__8_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_19__1__8_ccff_tail));

	tile_19__1_ tile_19__9_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[54:55]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[54:55]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[54:55]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__5_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__5_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_19__1__10_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__9_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__9_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_19__1__9_ccff_tail));

	tile_19__1_ tile_19__8_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[56:57]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[56:57]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[56:57]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__4_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__4_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_18__2__4_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__10_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__10_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_19__1__10_ccff_tail));

	tile_19__1_ tile_19__7_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[58:59]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[58:59]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[58:59]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__3_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__3_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_19__1__12_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__11_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__11_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_19__1__11_ccff_tail));

	tile_19__1_ tile_19__6_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[60:61]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[60:61]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[60:61]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__6__0_cby_18__6__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__6__0_cby_18__6__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_18__6__0_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__12_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__12_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_19__1__12_ccff_tail));

	tile_19__1_ tile_19__5_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[62:63]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[62:63]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[62:63]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_17__5__0_cby_18__5__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_17__5__0_cby_18__5__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_19__1__14_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__13_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__13_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(ccff_tail[8]));

	tile_19__1_ tile_19__4_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[64:65]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[64:65]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[64:65]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__2_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__2_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_18__2__2_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__14_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__14_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_19__1__14_ccff_tail));

	tile_19__1_ tile_19__3_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[66:67]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[66:67]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[66:67]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__1_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__1_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_19__1__16_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__15_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__15_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_19__1__15_ccff_tail));

	tile_19__1_ tile_19__2_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[68:69]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[68:69]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[68:69]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__0_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__0_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_18__2__0_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__16_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__16_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_19__1__16_ccff_tail));

	tile_19__1_ tile_19__1_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[70:71]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[70:71]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[70:71]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__1__0_cby_18__1__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__1__0_cby_18__1__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__0_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__17_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__17_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_19__1__17_ccff_tail));

	tile_1__0_ tile_18__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[72:73]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[72:73]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[72:73]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__1__0_cbx_18__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__1__0_cbx_18__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__1_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__0_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__0_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__0_ccff_tail));

	tile_1__0_ tile_17__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[74:75]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[74:75]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[74:75]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__16_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__16_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__2_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__1_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__1_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__1_ccff_tail));

	tile_1__0_ tile_16__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[76:77]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[76:77]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[76:77]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__15_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__15_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__3_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__2_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__2_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__2_ccff_tail));

	tile_1__0_ tile_15__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[78:79]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[78:79]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[78:79]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__14_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__14_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__4_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__3_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__3_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__3_ccff_tail));

	tile_1__0_ tile_14__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[80:81]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[80:81]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[80:81]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__13_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__13_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__5_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__4_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__4_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__4_ccff_tail));

	tile_1__0_ tile_13__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[82:83]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[82:83]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[82:83]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__12_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__12_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__6_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__5_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__5_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__5_ccff_tail));

	tile_1__0_ tile_12__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[84:85]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[84:85]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[84:85]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__11_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__11_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(ccff_head[1]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__6_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__6_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__6_ccff_tail));

	tile_1__0_ tile_11__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[86:87]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[86:87]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[86:87]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__10_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__10_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__8_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__7_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__7_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(ccff_tail[0]));

	tile_1__0_ tile_10__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[88:89]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[88:89]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[88:89]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__9_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__9_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__9_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__8_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__8_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__8_ccff_tail));

	tile_1__0_ tile_9__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[90:91]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[90:91]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[90:91]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__8_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__8_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__10_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__9_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__9_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__9_ccff_tail));

	tile_1__0_ tile_8__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[92:93]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[92:93]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[92:93]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__7_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__7_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__11_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__10_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__10_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__10_ccff_tail));

	tile_1__0_ tile_7__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[94:95]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[94:95]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[94:95]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__6_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__6_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__12_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__11_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__11_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__11_ccff_tail));

	tile_1__0_ tile_6__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[96:97]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[96:97]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[96:97]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__5_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__5_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__13_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__12_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__12_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__12_ccff_tail));

	tile_1__0_ tile_5__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[98:99]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[98:99]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[98:99]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__4_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__4_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__14_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__13_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__13_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__13_ccff_tail));

	tile_1__0_ tile_4__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[100:101]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[100:101]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[100:101]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__3_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__3_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__15_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__14_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__14_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__14_ccff_tail));

	tile_1__0_ tile_3__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[102:103]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[102:103]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[102:103]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__2_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__2_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__16_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__15_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__15_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__15_ccff_tail));

	tile_1__0_ tile_2__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[104:105]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[104:105]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[104:105]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__1_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__1_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__17_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__16_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__16_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__16_ccff_tail));

	tile_1__0_ tile_1__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[106:107]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[106:107]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[106:107]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__0_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__0_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(ccff_head[0]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__17_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__17_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__17_ccff_tail));

	tile_0__1_ tile_0__1_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[108:109]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[108:109]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[108:109]),
		.sb_0__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__17_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__17_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__0__chanx_right_in(tile_1__1__0_cbx_1__0__chanx_left_out[0:64]),
		.cby_0__1__chany_top_in(tile_0__2__0_sb_0__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__1__0_ccff_tail),
		.sb_0__0__chanx_right_out(tile_0__1__0_sb_0__0__chanx_right_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__1__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__1__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__1__chany_top_out(tile_0__1__0_cby_0__1__chany_top_out[0:64]),
		.ccff_tail(tile_0__1__0_ccff_tail));

	tile_0__2_ tile_0__2_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[110:111]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[110:111]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[110:111]),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__1__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__1__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__1__chanx_right_in(tile_1__2__0_cbx_1__1__chanx_left_out[0:64]),
		.sb_0__1__chany_bottom_in(tile_0__1__0_cby_0__1__chany_top_out[0:64]),
		.cby_0__2__chany_top_in(tile_0__2__1_sb_0__1__chany_bottom_out[0:64]),
		.ccff_head(tile_0__1__0_ccff_tail),
		.sb_0__1__chanx_right_out(tile_0__2__0_sb_0__1__chanx_right_out[0:64]),
		.sb_0__1__chany_bottom_out(tile_0__2__0_sb_0__1__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__2__chany_top_out(tile_0__2__0_cby_0__2__chany_top_out[0:64]),
		.ccff_tail(tile_0__2__0_ccff_tail));

	tile_0__2_ tile_0__3_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[112:113]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[112:113]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[112:113]),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__1__chanx_right_in(tile_1__2__1_cbx_1__1__chanx_left_out[0:64]),
		.sb_0__1__chany_bottom_in(tile_0__2__0_cby_0__2__chany_top_out[0:64]),
		.cby_0__2__chany_top_in(tile_0__2__2_sb_0__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[7]),
		.sb_0__1__chanx_right_out(tile_0__2__1_sb_0__1__chanx_right_out[0:64]),
		.sb_0__1__chany_bottom_out(tile_0__2__1_sb_0__1__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__1_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__1_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__2__chany_top_out(tile_0__2__1_cby_0__2__chany_top_out[0:64]),
		.ccff_tail(tile_0__2__1_ccff_tail));

	tile_0__2_ tile_0__4_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[114:115]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[114:115]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[114:115]),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__1_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__1_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__1__chanx_right_in(tile_1__2__2_cbx_1__1__chanx_left_out[0:64]),
		.sb_0__1__chany_bottom_in(tile_0__2__1_cby_0__2__chany_top_out[0:64]),
		.cby_0__2__chany_top_in(tile_0__5__0_sb_0__4__chany_bottom_out[0:64]),
		.ccff_head(tile_0__2__1_ccff_tail),
		.sb_0__1__chanx_right_out(tile_0__2__2_sb_0__1__chanx_right_out[0:64]),
		.sb_0__1__chany_bottom_out(tile_0__2__2_sb_0__1__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__2_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__2_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__2__chany_top_out(tile_0__2__2_cby_0__2__chany_top_out[0:64]),
		.ccff_tail(tile_0__2__2_ccff_tail));

	tile_0__2_ tile_0__7_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[120:121]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[120:121]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[120:121]),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__6__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__6__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__1__chanx_right_in(tile_1__2__3_cbx_1__1__chanx_left_out[0:64]),
		.sb_0__1__chany_bottom_in(tile_0__6__0_cby_0__6__chany_top_out[0:64]),
		.cby_0__2__chany_top_in(tile_0__2__4_sb_0__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__3_ccff_tail),
		.sb_0__1__chanx_right_out(tile_0__2__3_sb_0__1__chanx_right_out[0:64]),
		.sb_0__1__chany_bottom_out(tile_0__2__3_sb_0__1__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__3_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__3_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__2__chany_top_out(tile_0__2__3_cby_0__2__chany_top_out[0:64]),
		.ccff_tail(tile_0__2__3_ccff_tail));

	tile_0__2_ tile_0__8_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[122:123]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[122:123]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[122:123]),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__3_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__3_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__1__chanx_right_in(tile_1__2__4_cbx_1__1__chanx_left_out[0:64]),
		.sb_0__1__chany_bottom_in(tile_0__2__3_cby_0__2__chany_top_out[0:64]),
		.cby_0__2__chany_top_in(tile_0__2__5_sb_0__1__chany_bottom_out[0:64]),
		.ccff_head(tile_0__2__3_ccff_tail),
		.sb_0__1__chanx_right_out(tile_0__2__4_sb_0__1__chanx_right_out[0:64]),
		.sb_0__1__chany_bottom_out(tile_0__2__4_sb_0__1__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__4_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__4_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__2__chany_top_out(tile_0__2__4_cby_0__2__chany_top_out[0:64]),
		.ccff_tail(tile_0__2__4_ccff_tail));

	tile_0__2_ tile_0__9_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[124:125]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[124:125]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[124:125]),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__4_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__4_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__1__chanx_right_in(tile_1__2__5_cbx_1__1__chanx_left_out[0:64]),
		.sb_0__1__chany_bottom_in(tile_0__2__4_cby_0__2__chany_top_out[0:64]),
		.cby_0__2__chany_top_in(tile_0__10__0_sb_0__9__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__5_ccff_tail),
		.sb_0__1__chanx_right_out(tile_0__2__5_sb_0__1__chanx_right_out[0:64]),
		.sb_0__1__chany_bottom_out(tile_0__2__5_sb_0__1__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__5_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__5_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__2__chany_top_out(tile_0__2__5_cby_0__2__chany_top_out[0:64]),
		.ccff_tail(tile_0__2__5_ccff_tail));

	tile_0__2_ tile_0__12_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[130:131]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[130:131]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[130:131]),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__11__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__11__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__1__chanx_right_in(tile_1__2__6_cbx_1__1__chanx_left_out[0:64]),
		.sb_0__1__chany_bottom_in(tile_0__11__0_cby_0__11__chany_top_out[0:64]),
		.cby_0__2__chany_top_in(tile_0__2__7_sb_0__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[20]),
		.sb_0__1__chanx_right_out(tile_0__2__6_sb_0__1__chanx_right_out[0:64]),
		.sb_0__1__chany_bottom_out(tile_0__2__6_sb_0__1__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__6_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__6_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__2__chany_top_out(tile_0__2__6_cby_0__2__chany_top_out[0:64]),
		.ccff_tail(tile_0__2__6_ccff_tail));

	tile_0__2_ tile_0__13_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[132:133]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[132:133]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[132:133]),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__6_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__6_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__1__chanx_right_in(tile_1__2__7_cbx_1__1__chanx_left_out[0:64]),
		.sb_0__1__chany_bottom_in(tile_0__2__6_cby_0__2__chany_top_out[0:64]),
		.cby_0__2__chany_top_in(tile_0__5__1_sb_0__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__7_ccff_tail),
		.sb_0__1__chanx_right_out(tile_0__2__7_sb_0__1__chanx_right_out[0:64]),
		.sb_0__1__chany_bottom_out(tile_0__2__7_sb_0__1__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__7_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__7_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__2__chany_top_out(tile_0__2__7_cby_0__2__chany_top_out[0:64]),
		.ccff_tail(tile_0__2__7_ccff_tail));

	tile_0__2_ tile_0__16_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[138:139]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[138:139]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[138:139]),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__6__1_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__6__1_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__1__chanx_right_in(tile_1__2__8_cbx_1__1__chanx_left_out[0:64]),
		.sb_0__1__chany_bottom_in(tile_0__6__1_cby_0__6__chany_top_out[0:64]),
		.cby_0__2__chany_top_in(tile_0__2__9_sb_0__1__chany_bottom_out[0:64]),
		.ccff_head(tile_0__6__1_ccff_tail),
		.sb_0__1__chanx_right_out(tile_0__2__8_sb_0__1__chanx_right_out[0:64]),
		.sb_0__1__chany_bottom_out(tile_0__2__8_sb_0__1__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__8_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__8_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__2__chany_top_out(tile_0__2__8_cby_0__2__chany_top_out[0:64]),
		.ccff_tail(tile_0__2__8_ccff_tail));

	tile_0__2_ tile_0__17_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[140:141]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[140:141]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[140:141]),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__8_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__8_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__1__chanx_right_in(tile_1__2__9_cbx_1__1__chanx_left_out[0:64]),
		.sb_0__1__chany_bottom_in(tile_0__2__8_cby_0__2__chany_top_out[0:64]),
		.cby_0__2__chany_top_in(tile_0__2__10_sb_0__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[30]),
		.sb_0__1__chanx_right_out(tile_0__2__9_sb_0__1__chanx_right_out[0:64]),
		.sb_0__1__chany_bottom_out(tile_0__2__9_sb_0__1__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__9_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__9_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__2__chany_top_out(tile_0__2__9_cby_0__2__chany_top_out[0:64]),
		.ccff_tail(tile_0__2__9_ccff_tail));

	tile_0__2_ tile_0__18_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[142:143]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[142:143]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[142:143]),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__9_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__9_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__1__chanx_right_in(tile_1__2__10_cbx_1__1__chanx_left_out[0:64]),
		.sb_0__1__chany_bottom_in(tile_0__2__9_cby_0__2__chany_top_out[0:64]),
		.cby_0__2__chany_top_in(tile_0__19__0_sb_0__18__chany_bottom_out[0:64]),
		.ccff_head(tile_0__2__9_ccff_tail),
		.sb_0__1__chanx_right_out(tile_0__2__10_sb_0__1__chanx_right_out[0:64]),
		.sb_0__1__chany_bottom_out(tile_0__2__10_sb_0__1__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__10_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__10_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__2__chany_top_out(tile_0__2__10_cby_0__2__chany_top_out[0:64]),
		.ccff_tail(tile_0__2__10_ccff_tail));

	tile_0__5_ tile_0__5_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[116:117]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[116:117]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[116:117]),
		.sb_0__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__2_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__4__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__2_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__4__chanx_right_in(tile_1__5__0_cbx_1__4__chanx_left_out[0:64]),
		.sb_0__4__chany_bottom_in(tile_0__2__2_cby_0__2__chany_top_out[0:64]),
		.cby_0__5__chany_top_in(tile_0__6__0_sb_0__5__chany_bottom_out[0:64]),
		.ccff_head(tile_1__5__0_ccff_tail),
		.sb_0__4__chanx_right_out(tile_0__5__0_sb_0__4__chanx_right_out[0:64]),
		.sb_0__4__chany_bottom_out(tile_0__5__0_sb_0__4__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__5__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__5__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__5__chany_top_out(tile_0__5__0_cby_0__5__chany_top_out[0:64]),
		.ccff_tail(tile_0__5__0_ccff_tail));

	tile_0__5_ tile_0__14_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[134:135]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[134:135]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[134:135]),
		.sb_0__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__7_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__4__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__7_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__4__chanx_right_in(tile_1__5__1_cbx_1__4__chanx_left_out[0:64]),
		.sb_0__4__chany_bottom_in(tile_0__2__7_cby_0__2__chany_top_out[0:64]),
		.cby_0__5__chany_top_in(tile_0__6__1_sb_0__5__chany_bottom_out[0:64]),
		.ccff_head(tile_0__2__7_ccff_tail),
		.sb_0__4__chanx_right_out(tile_0__5__1_sb_0__4__chanx_right_out[0:64]),
		.sb_0__4__chany_bottom_out(tile_0__5__1_sb_0__4__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__5__1_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__5__1_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__5__chany_top_out(tile_0__5__1_cby_0__5__chany_top_out[0:64]),
		.ccff_tail(tile_0__5__1_ccff_tail));

	tile_0__6_ tile_0__6_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[118:119]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[118:119]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[118:119]),
		.sb_0__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_0__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_0__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_0__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_0__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_0__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_0__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_0__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_0__5__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__5__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__5__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__5__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__5__chanx_right_in(tile_1__6__0_cbx_1__5__chanx_left_out[0:64]),
		.sb_0__5__chany_bottom_in(tile_0__5__0_cby_0__5__chany_top_out[0:64]),
		.cby_0__6__chany_top_in(tile_0__2__3_sb_0__1__chany_bottom_out[0:64]),
		.ccff_head(tile_0__5__0_ccff_tail),
		.sb_0__5__chanx_right_out(tile_0__6__0_sb_0__5__chanx_right_out[0:64]),
		.sb_0__5__chany_bottom_out(tile_0__6__0_sb_0__5__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__6__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__6__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__6__chany_top_out(tile_0__6__0_cby_0__6__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[9]));

	tile_0__6_ tile_0__15_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[136:137]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[136:137]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[136:137]),
		.sb_0__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_0__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_0__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_0__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_0__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_0__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_0__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_0__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_0__5__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__5__1_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__5__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__5__1_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__5__chanx_right_in(tile_1__6__1_cbx_1__5__chanx_left_out[0:64]),
		.sb_0__5__chany_bottom_in(tile_0__5__1_cby_0__5__chany_top_out[0:64]),
		.cby_0__6__chany_top_in(tile_0__2__8_sb_0__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__6__1_ccff_tail),
		.sb_0__5__chanx_right_out(tile_0__6__1_sb_0__5__chanx_right_out[0:64]),
		.sb_0__5__chany_bottom_out(tile_0__6__1_sb_0__5__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__6__1_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__6__1_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__6__chany_top_out(tile_0__6__1_cby_0__6__chany_top_out[0:64]),
		.ccff_tail(tile_0__6__1_ccff_tail));

	tile_0__10_ tile_0__10_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[126:127]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[126:127]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[126:127]),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.sb_0__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.sb_0__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__5_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__9__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__5_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__9__chanx_right_in(tile_1__10__0_cbx_1__9__chanx_left_out[0:64]),
		.sb_0__9__chany_bottom_in(tile_0__2__5_cby_0__2__chany_top_out[0:64]),
		.cby_0__10__chany_top_in(tile_0__11__0_sb_0__10__chany_bottom_out[0:64]),
		.ccff_head(tile_0__2__5_ccff_tail),
		.sb_0__9__chanx_right_out(tile_0__10__0_sb_0__9__chanx_right_out[0:64]),
		.sb_0__9__chany_bottom_out(tile_0__10__0_sb_0__9__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__10__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__10__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__10__chany_top_out(tile_0__10__0_cby_0__10__chany_top_out[0:64]),
		.ccff_tail(tile_0__10__0_ccff_tail));

	tile_0__11_ tile_0__11_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[128:129]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[128:129]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[128:129]),
		.sb_0__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__10__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__10__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__10__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__10__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__10__chanx_right_in(tile_1__11__0_cbx_1__10__chanx_left_out[0:64]),
		.sb_0__10__chany_bottom_in(tile_0__10__0_cby_0__10__chany_top_out[0:64]),
		.cby_0__11__chany_top_in(tile_0__2__6_sb_0__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__11__0_ccff_tail),
		.sb_0__10__chanx_right_out(tile_0__11__0_sb_0__10__chanx_right_out[0:64]),
		.sb_0__10__chany_bottom_out(tile_0__11__0_sb_0__10__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__11__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__11__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__11__chany_top_out(tile_0__11__0_cby_0__11__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[19]));

	tile_1__1_ tile_1__1_ (
		.prog_clk(prog_clk),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__16_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__16_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__17_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__17_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__chanx_right_in(tile_1__1__1_cbx_1__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_0_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__0__chanx_left_in(tile_0__1__0_sb_0__0__chanx_right_out[0:64]),
		.cby_1__1__chany_top_in(tile_1__2__0_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__1__1_ccff_tail),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__0_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__0_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_1__0__chanx_right_out(tile_1__1__0_sb_1__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__0__chanx_left_out(tile_1__1__0_cbx_1__0__chanx_left_out[0:64]),
		.cby_1__1__chany_top_out(tile_1__1__0_cby_1__1__chany_top_out[0:64]),
		.ccff_tail(tile_1__1__0_ccff_tail));

	tile_1__1_ tile_2__1_ (
		.prog_clk(prog_clk),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__15_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__15_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__16_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__16_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__chanx_right_in(tile_1__1__2_cbx_1__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_11_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__0__chanx_left_in(tile_1__1__0_sb_1__0__chanx_right_out[0:64]),
		.cby_1__1__chany_top_in(tile_1__2__11_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__1__2_ccff_tail),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__1_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__1_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_1__0__chanx_right_out(tile_1__1__1_sb_1__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_2__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__0__chanx_left_out(tile_1__1__1_cbx_1__0__chanx_left_out[0:64]),
		.cby_1__1__chany_top_out(tile_1__1__1_cby_1__1__chany_top_out[0:64]),
		.ccff_tail(tile_1__1__1_ccff_tail));

	tile_1__1_ tile_3__1_ (
		.prog_clk(prog_clk),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__14_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__14_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__15_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__15_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__chanx_right_in(tile_1__1__3_cbx_1__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_22_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__0__chanx_left_in(tile_1__1__1_sb_1__0__chanx_right_out[0:64]),
		.cby_1__1__chany_top_in(tile_1__2__22_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__1__3_ccff_tail),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__2_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__2_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_1__0__chanx_right_out(tile_1__1__2_sb_1__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_3__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__0__chanx_left_out(tile_1__1__2_cbx_1__0__chanx_left_out[0:64]),
		.cby_1__1__chany_top_out(tile_1__1__2_cby_1__1__chany_top_out[0:64]),
		.ccff_tail(tile_1__1__2_ccff_tail));

	tile_1__1_ tile_4__1_ (
		.prog_clk(prog_clk),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__13_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__13_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__14_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__14_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__chanx_right_in(tile_1__1__4_cbx_1__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_33_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__0__chanx_left_in(tile_1__1__2_sb_1__0__chanx_right_out[0:64]),
		.cby_1__1__chany_top_in(tile_1__2__33_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[3]),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__3_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__3_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_1__0__chanx_right_out(tile_1__1__3_sb_1__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_4__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__0__chanx_left_out(tile_1__1__3_cbx_1__0__chanx_left_out[0:64]),
		.cby_1__1__chany_top_out(tile_1__1__3_cby_1__1__chany_top_out[0:64]),
		.ccff_tail(tile_1__1__3_ccff_tail));

	tile_1__1_ tile_5__1_ (
		.prog_clk(prog_clk),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__12_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__12_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__13_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__13_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__chanx_right_in(tile_1__1__5_cbx_1__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_44_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__0__chanx_left_in(tile_1__1__3_sb_1__0__chanx_right_out[0:64]),
		.cby_1__1__chany_top_in(tile_1__2__44_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__1__5_ccff_tail),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__4_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__4_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_1__0__chanx_right_out(tile_1__1__4_sb_1__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_5__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__0__chanx_left_out(tile_1__1__4_cbx_1__0__chanx_left_out[0:64]),
		.cby_1__1__chany_top_out(tile_1__1__4_cby_1__1__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[2]));

	tile_1__1_ tile_6__1_ (
		.prog_clk(prog_clk),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__11_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__11_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__12_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__12_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__chanx_right_in(tile_1__1__6_cbx_1__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_55_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__0__chanx_left_in(tile_1__1__4_sb_1__0__chanx_right_out[0:64]),
		.cby_1__1__chany_top_in(tile_1__2__55_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__1__6_ccff_tail),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__5_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__5_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_1__0__chanx_right_out(tile_1__1__5_sb_1__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_6__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__0__chanx_left_out(tile_1__1__5_cbx_1__0__chanx_left_out[0:64]),
		.cby_1__1__chany_top_out(tile_1__1__5_cby_1__1__chany_top_out[0:64]),
		.ccff_tail(tile_1__1__5_ccff_tail));

	tile_1__1_ tile_7__1_ (
		.prog_clk(prog_clk),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__10_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__10_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__11_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__11_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__chanx_right_in(tile_1__1__7_cbx_1__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_66_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__0__chanx_left_in(tile_1__1__5_sb_1__0__chanx_right_out[0:64]),
		.cby_1__1__chany_top_in(tile_1__2__66_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__1__7_ccff_tail),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__6_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__6_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_1__0__chanx_right_out(tile_1__1__6_sb_1__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_7__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__0__chanx_left_out(tile_1__1__6_cbx_1__0__chanx_left_out[0:64]),
		.cby_1__1__chany_top_out(tile_1__1__6_cby_1__1__chany_top_out[0:64]),
		.ccff_tail(tile_1__1__6_ccff_tail));

	tile_1__1_ tile_8__1_ (
		.prog_clk(prog_clk),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__9_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__9_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__10_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__10_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__chanx_right_in(tile_1__1__8_cbx_1__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_77_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__0__chanx_left_in(tile_1__1__6_sb_1__0__chanx_right_out[0:64]),
		.cby_1__1__chany_top_in(tile_1__2__77_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__1__8_ccff_tail),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__7_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__7_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_1__0__chanx_right_out(tile_1__1__7_sb_1__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_8__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__0__chanx_left_out(tile_1__1__7_cbx_1__0__chanx_left_out[0:64]),
		.cby_1__1__chany_top_out(tile_1__1__7_cby_1__1__chany_top_out[0:64]),
		.ccff_tail(tile_1__1__7_ccff_tail));

	tile_1__1_ tile_9__1_ (
		.prog_clk(prog_clk),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__8_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__8_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__9_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__9_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__chanx_right_in(tile_1__1__9_cbx_1__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_88_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__0__chanx_left_in(tile_1__1__7_sb_1__0__chanx_right_out[0:64]),
		.cby_1__1__chany_top_in(tile_1__2__88_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__1__9_ccff_tail),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__8_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__8_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_1__0__chanx_right_out(tile_1__1__8_sb_1__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_9__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__0__chanx_left_out(tile_1__1__8_cbx_1__0__chanx_left_out[0:64]),
		.cby_1__1__chany_top_out(tile_1__1__8_cby_1__1__chany_top_out[0:64]),
		.ccff_tail(tile_1__1__8_ccff_tail));

	tile_1__1_ tile_10__1_ (
		.prog_clk(prog_clk),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__7_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__7_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__8_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__8_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__chanx_right_in(tile_1__1__10_cbx_1__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_99_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__0__chanx_left_in(tile_1__1__8_sb_1__0__chanx_right_out[0:64]),
		.cby_1__1__chany_top_in(tile_1__2__99_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__1__10_ccff_tail),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__9_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__9_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_1__0__chanx_right_out(tile_1__1__9_sb_1__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_10__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__0__chanx_left_out(tile_1__1__9_cbx_1__0__chanx_left_out[0:64]),
		.cby_1__1__chany_top_out(tile_1__1__9_cby_1__1__chany_top_out[0:64]),
		.ccff_tail(tile_1__1__9_ccff_tail));

	tile_1__1_ tile_11__1_ (
		.prog_clk(prog_clk),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__6_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__6_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__7_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__7_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__chanx_right_in(tile_1__1__11_cbx_1__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_110_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__0__chanx_left_in(tile_1__1__9_sb_1__0__chanx_right_out[0:64]),
		.cby_1__1__chany_top_in(tile_1__2__110_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__1__11_ccff_tail),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__10_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__10_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_1__0__chanx_right_out(tile_1__1__10_sb_1__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_11__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__0__chanx_left_out(tile_1__1__10_cbx_1__0__chanx_left_out[0:64]),
		.cby_1__1__chany_top_out(tile_1__1__10_cby_1__1__chany_top_out[0:64]),
		.ccff_tail(tile_1__1__10_ccff_tail));

	tile_1__1_ tile_12__1_ (
		.prog_clk(prog_clk),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__5_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__5_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__6_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__6_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__chanx_right_in(tile_1__1__12_cbx_1__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_121_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__0__chanx_left_in(tile_1__1__10_sb_1__0__chanx_right_out[0:64]),
		.cby_1__1__chany_top_in(tile_1__2__121_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__1__12_ccff_tail),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__11_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__11_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_1__0__chanx_right_out(tile_1__1__11_sb_1__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_12__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__0__chanx_left_out(tile_1__1__11_cbx_1__0__chanx_left_out[0:64]),
		.cby_1__1__chany_top_out(tile_1__1__11_cby_1__1__chany_top_out[0:64]),
		.ccff_tail(tile_1__1__11_ccff_tail));

	tile_1__1_ tile_13__1_ (
		.prog_clk(prog_clk),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__4_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__4_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__5_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__5_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__chanx_right_in(tile_1__1__13_cbx_1__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_132_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__0__chanx_left_in(tile_1__1__11_sb_1__0__chanx_right_out[0:64]),
		.cby_1__1__chany_top_in(tile_1__2__132_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__1__13_ccff_tail),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__12_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__12_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_1__0__chanx_right_out(tile_1__1__12_sb_1__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_13__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__0__chanx_left_out(tile_1__1__12_cbx_1__0__chanx_left_out[0:64]),
		.cby_1__1__chany_top_out(tile_1__1__12_cby_1__1__chany_top_out[0:64]),
		.ccff_tail(tile_1__1__12_ccff_tail));

	tile_1__1_ tile_14__1_ (
		.prog_clk(prog_clk),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__3_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__3_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__4_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__4_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__chanx_right_in(tile_1__1__14_cbx_1__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_143_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__0__chanx_left_in(tile_1__1__12_sb_1__0__chanx_right_out[0:64]),
		.cby_1__1__chany_top_in(tile_1__2__143_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__1__14_ccff_tail),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__13_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__13_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_1__0__chanx_right_out(tile_1__1__13_sb_1__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_14__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__0__chanx_left_out(tile_1__1__13_cbx_1__0__chanx_left_out[0:64]),
		.cby_1__1__chany_top_out(tile_1__1__13_cby_1__1__chany_top_out[0:64]),
		.ccff_tail(tile_1__1__13_ccff_tail));

	tile_1__1_ tile_15__1_ (
		.prog_clk(prog_clk),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__2_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__2_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__3_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__3_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__chanx_right_in(tile_1__1__15_cbx_1__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_154_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__0__chanx_left_in(tile_1__1__13_sb_1__0__chanx_right_out[0:64]),
		.cby_1__1__chany_top_in(tile_1__2__154_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[2]),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__14_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__14_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_1__0__chanx_right_out(tile_1__1__14_sb_1__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_15__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__0__chanx_left_out(tile_1__1__14_cbx_1__0__chanx_left_out[0:64]),
		.cby_1__1__chany_top_out(tile_1__1__14_cby_1__1__chany_top_out[0:64]),
		.ccff_tail(tile_1__1__14_ccff_tail));

	tile_1__1_ tile_16__1_ (
		.prog_clk(prog_clk),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__1_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__1_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__2_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__2_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__chanx_right_in(tile_1__1__16_cbx_1__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_165_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__0__chanx_left_in(tile_1__1__14_sb_1__0__chanx_right_out[0:64]),
		.cby_1__1__chany_top_in(tile_1__2__165_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__1__16_ccff_tail),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__15_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__15_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_1__0__chanx_right_out(tile_1__1__15_sb_1__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_16__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__0__chanx_left_out(tile_1__1__15_cbx_1__0__chanx_left_out[0:64]),
		.cby_1__1__chany_top_out(tile_1__1__15_cby_1__1__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[1]));

	tile_1__1_ tile_17__1_ (
		.prog_clk(prog_clk),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__0_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__0_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__1_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__1_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__chanx_right_in(tile_18__1__0_cbx_18__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_176_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__0__chanx_left_in(tile_1__1__15_sb_1__0__chanx_right_out[0:64]),
		.cby_1__1__chany_top_in(tile_1__2__176_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_18__1__0_ccff_tail),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__16_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__16_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_1__0__chanx_right_out(tile_1__1__16_sb_1__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_17__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__0__chanx_left_out(tile_1__1__16_cbx_1__0__chanx_left_out[0:64]),
		.cby_1__1__chany_top_out(tile_1__1__16_cby_1__1__chany_top_out[0:64]),
		.ccff_tail(tile_1__1__16_ccff_tail));

	tile_1__2_ tile_1__2_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__11_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__1__0_cby_1__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_1_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_0__2__0_sb_0__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__1_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_0__2__0_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__0_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__0_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__0_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__0_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__0_ccff_tail));

	tile_1__2_ tile_1__3_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__12_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__0_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_2_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_0__2__1_sb_0__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__2_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__12_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__1_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__1_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__1_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__1_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[6]));

	tile_1__2_ tile_1__4_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__13_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__1_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_1__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_0__2__2_sb_0__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__0_sb_1__4__chany_bottom_out[0:64]),
		.ccff_head(tile_0__2__2_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__2_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__2_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__2_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__2_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__2_ccff_tail));

	tile_1__2_ tile_1__7_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__14_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__6__0_cby_1__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_4_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_0__2__3_sb_0__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__4_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__14_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__3_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__3_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__3_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__3_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__3_ccff_tail));

	tile_1__2_ tile_1__8_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__15_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__3_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_5_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_0__2__4_sb_0__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__5_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_0__2__4_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__4_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__4_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__4_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__4_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__4_ccff_tail));

	tile_1__2_ tile_1__9_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__16_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__4_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_1__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_0__2__5_sb_0__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__10__0_sb_1__9__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[17]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__5_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__5_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__5_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__5_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__5_ccff_tail));

	tile_1__2_ tile_1__12_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__17_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__11__0_cby_1__11__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_7_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_0__2__6_sb_0__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__7_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_0__2__6_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__6_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__6_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__6_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__6_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__6_ccff_tail));

	tile_1__2_ tile_1__13_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__18_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__18_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__18_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__18_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__18_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__18_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__18_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__6_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_1__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_0__2__7_sb_0__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__1_sb_1__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__18_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__7_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__7_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__7_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__7_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__7_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__7_ccff_tail));

	tile_1__2_ tile_1__16_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__19_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__19_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__19_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__19_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__19_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__19_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__19_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__6__1_cby_1__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_9_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_0__2__8_sb_0__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__9_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_0__2__8_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__8_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__8_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__8_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__8_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__8_ccff_tail));

	tile_1__2_ tile_1__17_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__20_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__20_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__20_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__20_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__20_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__20_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__20_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__8_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_10_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_0__2__9_sb_0__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__10_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__20_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__9_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__9_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__9_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__9_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__9_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[29]));

	tile_1__2_ tile_1__18_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__21_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__21_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__21_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__21_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__21_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__21_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__21_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__9_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__0_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_1__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_0__2__10_sb_0__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__19__0_sb_1__18__chany_bottom_out[0:64]),
		.ccff_head(tile_0__2__10_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__10_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__10_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__10_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__10_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__10_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__10_ccff_tail));

	tile_1__2_ tile_2__2_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__22_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__22_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__22_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__22_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__22_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__22_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__22_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__1__1_cby_1__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_12_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__0_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__12_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__0_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__11_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__11_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__11_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__11_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__11_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__11_ccff_tail));

	tile_1__2_ tile_2__3_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__23_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__23_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__23_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__23_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__23_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__23_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__23_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__11_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_13_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__1_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__13_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__23_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__12_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__12_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__12_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__12_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__12_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__12_ccff_tail));

	tile_1__2_ tile_2__4_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__24_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__24_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__24_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__24_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__24_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__24_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__24_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__12_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_2__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__2_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__0_sb_2__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__2_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__13_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__13_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__13_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__13_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__13_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__13_ccff_tail));

	tile_1__2_ tile_2__7_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__25_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__25_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__25_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__25_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__25_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__25_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__25_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__6__0_cby_2__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_15_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__3_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__15_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__25_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__14_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__14_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__14_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__14_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__14_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__14_ccff_tail));

	tile_1__2_ tile_2__8_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__26_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__26_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__26_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__26_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__26_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__26_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__26_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__14_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_16_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__4_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__16_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__4_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__15_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__15_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__15_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__15_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__15_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__15_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__15_ccff_tail));

	tile_1__2_ tile_2__9_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__27_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__27_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__27_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__27_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__27_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__27_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__27_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__15_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_2__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__5_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__10__0_sb_2__9__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__27_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__16_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__16_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__16_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__16_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__16_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__16_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[16]));

	tile_1__2_ tile_2__12_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__28_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__28_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__28_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__28_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__28_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__28_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__28_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__11__0_cby_2__11__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_18_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__6_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__18_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__6_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__17_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__17_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__17_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__17_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__17_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__17_ccff_tail));

	tile_1__2_ tile_2__13_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__29_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__29_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__29_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__29_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__29_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__29_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__29_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__17_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_2__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__7_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__1_sb_2__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__29_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__18_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__18_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__18_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__18_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__18_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__18_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__18_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__18_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__18_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__18_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__18_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__18_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__18_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__18_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__18_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__18_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__18_ccff_tail));

	tile_1__2_ tile_2__16_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__30_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__30_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__30_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__30_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__30_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__30_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__30_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__6__1_cby_2__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_20_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__8_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__20_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__8_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__19_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__19_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__19_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__19_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__19_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__19_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__19_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__19_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__19_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__19_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__19_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__19_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__19_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__19_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__19_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__19_ccff_tail));

	tile_1__2_ tile_2__17_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__31_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__31_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__31_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__31_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__31_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__31_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__19_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__19_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__19_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__19_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__19_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__31_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__19_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_21_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__9_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__21_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__31_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__20_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__20_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__20_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__20_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__20_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__20_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__20_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__20_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__20_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__20_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__20_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__20_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__20_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__20_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__20_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__20_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__20_ccff_tail));

	tile_1__2_ tile_2__18_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__32_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__32_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__32_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__32_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__32_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__32_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__20_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__20_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__20_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__20_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__20_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__32_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__20_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__1_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_2__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__10_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__19__1_sb_1__18__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__10_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__21_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__21_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__21_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__21_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__21_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__21_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__21_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__21_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__21_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__21_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__21_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__21_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__21_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__21_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__21_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__21_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__21_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__21_ccff_tail));

	tile_1__2_ tile_3__2_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__33_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__33_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__33_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__33_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__33_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__33_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__33_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__1__2_cby_1__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_23_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__11_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__23_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__11_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__22_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__22_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__22_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__22_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__22_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__22_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__22_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__22_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__22_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__22_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__22_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__22_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__22_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__22_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__22_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__22_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__22_ccff_tail));

	tile_1__2_ tile_3__3_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__34_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__34_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__34_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__34_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__34_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__34_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__22_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__22_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__22_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__22_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__22_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__34_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__22_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_24_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__12_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__24_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__34_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__23_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__23_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__23_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__23_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__23_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__23_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__23_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__23_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__23_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__23_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__23_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__23_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__23_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__23_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__23_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__23_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__23_ccff_tail));

	tile_1__2_ tile_3__4_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__35_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__35_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__35_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__35_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__35_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__35_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__23_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__23_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__23_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__23_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__23_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__35_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__23_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_3__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__13_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__2_sb_1__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__13_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__24_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__24_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__24_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__24_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__24_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__24_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__24_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__24_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__24_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__24_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__24_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__24_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__24_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__24_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__24_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__24_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__24_ccff_tail));

	tile_1__2_ tile_3__7_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__36_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__36_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__36_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__36_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__36_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__36_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__36_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__6__2_cby_1__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_26_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__14_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__26_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__36_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__25_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__25_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__25_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__25_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__25_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__25_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__25_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__25_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__25_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__25_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__25_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__25_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__25_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__25_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__25_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__25_ccff_tail));

	tile_1__2_ tile_3__8_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__37_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__37_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__37_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__37_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__37_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__37_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__25_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__25_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__25_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__25_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__25_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__37_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__25_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_27_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__15_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__27_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__15_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__26_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__26_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__26_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__26_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__26_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__26_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__26_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__26_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__26_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__26_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__26_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__26_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__26_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__26_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__26_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__26_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__26_ccff_tail));

	tile_1__2_ tile_3__9_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__38_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__38_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__38_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__38_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__38_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__38_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__26_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__26_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__26_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__26_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__26_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__38_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__26_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_3__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__16_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__10__1_sb_1__9__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__38_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__27_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__27_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__27_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__27_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__27_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__27_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__27_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__27_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__27_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__27_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__27_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__27_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__27_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__27_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__27_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__27_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__27_ccff_tail));

	tile_1__2_ tile_3__12_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__39_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__39_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__39_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__39_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__39_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__39_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__39_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__11__1_cby_1__11__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_29_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__17_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__29_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__17_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__28_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__28_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__28_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__28_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__28_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__28_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__28_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__28_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__28_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__28_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__28_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__28_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__28_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__28_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__28_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__28_ccff_tail));

	tile_1__2_ tile_3__13_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__40_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__40_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__40_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__40_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__40_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__40_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__28_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__28_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__28_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__28_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__28_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__40_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__28_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_3__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__18_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__3_sb_1__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__40_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__29_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__29_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__29_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__29_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__29_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__29_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__29_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__29_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__29_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__29_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__29_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__29_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__29_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__29_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__29_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__29_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__29_ccff_tail));

	tile_1__2_ tile_3__16_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__41_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__41_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__41_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__41_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__41_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__41_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__41_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__6__3_cby_1__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_31_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__19_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__31_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__19_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__30_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__30_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__30_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__30_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__30_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__30_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__30_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__30_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__30_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__30_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__30_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__30_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__30_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__30_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__30_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__30_ccff_tail));

	tile_1__2_ tile_3__17_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__42_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__42_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__42_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__42_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__42_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__42_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__30_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__30_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__30_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__30_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__30_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__42_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__30_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_32_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__20_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__32_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__42_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__31_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__31_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__31_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__31_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__31_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__31_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__31_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__31_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__31_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__31_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__31_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__31_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__31_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__31_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__31_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__31_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__31_ccff_tail));

	tile_1__2_ tile_3__18_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__43_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__43_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__43_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__43_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__43_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__43_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__31_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__31_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__31_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__31_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__31_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__43_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__31_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__2_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_3__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__21_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__19__2_sb_1__18__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__21_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__32_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__32_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__32_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__32_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__32_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__32_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__32_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__32_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__32_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__32_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__32_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__32_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__32_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__32_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__32_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__32_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__32_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__32_ccff_tail));

	tile_1__2_ tile_4__2_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__44_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__44_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__44_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__44_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__44_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__44_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__44_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__1__3_cby_1__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_34_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__22_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__34_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__22_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__33_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__33_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__33_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__33_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__33_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__33_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__33_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__33_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__33_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__33_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__33_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__33_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__33_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__33_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__33_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__33_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__33_ccff_tail));

	tile_1__2_ tile_4__3_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__45_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__45_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__45_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__45_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__45_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__45_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__33_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__33_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__33_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__33_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__33_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__45_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__33_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_35_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__23_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__35_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__45_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__34_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__34_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__34_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__34_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__34_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__34_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__34_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__34_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__34_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__34_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__34_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__34_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__34_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__34_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__34_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__34_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__34_ccff_tail));

	tile_1__2_ tile_4__4_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__46_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__46_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__46_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__46_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__46_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__46_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__34_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__34_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__34_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__34_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__34_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__46_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__34_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_4__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__24_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__2_sb_2__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__24_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__35_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__35_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__35_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__35_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__35_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__35_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__35_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__35_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__35_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__35_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__35_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__35_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__35_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__35_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__35_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__35_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__35_ccff_tail));

	tile_1__2_ tile_4__7_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__47_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__47_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__47_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__47_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__47_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__47_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__47_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__6__2_cby_2__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_37_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__25_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__37_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__47_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__36_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__36_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__36_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__36_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__36_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__36_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__36_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__36_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__36_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__36_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__36_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__36_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__36_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__36_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__36_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__36_ccff_tail));

	tile_1__2_ tile_4__8_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__48_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__48_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__48_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__48_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__48_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__48_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__36_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__36_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__36_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__36_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__36_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__48_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__36_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_38_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__26_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__38_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__26_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__37_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__37_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__37_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__37_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__37_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__37_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__37_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__37_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__37_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__37_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__37_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__37_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__37_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__37_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__37_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__37_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[13]));

	tile_1__2_ tile_4__9_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__49_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__49_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__49_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__49_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__49_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__49_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__37_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__37_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__37_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__37_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__37_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__49_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__37_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_4__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__27_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__10__1_sb_2__9__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__49_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__38_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__38_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__38_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__38_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__38_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__38_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__38_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__38_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__38_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__38_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__38_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__38_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__38_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__38_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__38_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__38_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__38_ccff_tail));

	tile_1__2_ tile_4__12_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__50_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__50_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__50_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__50_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__50_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__50_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__50_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__11__1_cby_2__11__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_40_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__28_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__40_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__28_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__39_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__39_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__39_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__39_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__39_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__39_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__39_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__39_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__39_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__39_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__39_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__39_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__39_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__39_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__39_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__39_ccff_tail));

	tile_1__2_ tile_4__13_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__51_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__51_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__51_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__51_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__51_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__51_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__39_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__39_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__39_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__39_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__39_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__51_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__39_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_4__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__29_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__3_sb_2__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__51_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__40_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__40_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__40_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__40_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__40_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__40_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__40_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__40_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__40_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__40_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__40_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__40_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__40_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__40_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__40_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__40_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__40_ccff_tail));

	tile_1__2_ tile_4__16_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__52_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__52_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__52_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__52_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__52_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__52_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__52_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__6__3_cby_2__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_42_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__30_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__42_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__30_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__41_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__41_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__41_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__41_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__41_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__41_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__41_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__41_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__41_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__41_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__41_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__41_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__41_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__41_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__41_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__41_ccff_tail));

	tile_1__2_ tile_4__17_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__53_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__53_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__53_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__53_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__53_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__53_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__41_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__41_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__41_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__41_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__41_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__53_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__41_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_43_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__31_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__43_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__53_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__42_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__42_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__42_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__42_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__42_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__42_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__42_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__42_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__42_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__42_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__42_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__42_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__42_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__42_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__42_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__42_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__42_ccff_tail));

	tile_1__2_ tile_4__18_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__54_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__54_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__54_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__54_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__54_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__54_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__42_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__42_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__42_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__42_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__42_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__54_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__42_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__3_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_4__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__32_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__19__3_sb_1__18__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__32_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__43_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__43_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__43_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__43_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__43_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__43_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__43_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__43_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__43_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__43_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__43_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__43_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__43_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__43_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__43_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__43_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__43_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__43_ccff_tail));

	tile_1__2_ tile_5__2_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__55_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__55_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__55_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__55_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__55_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__55_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__55_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__1__4_cby_1__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_45_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__33_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__45_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__33_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__44_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__44_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__44_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__44_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__44_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__44_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__44_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__44_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__44_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__44_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__44_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__44_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__44_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__44_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__44_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__44_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[3]));

	tile_1__2_ tile_5__3_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__56_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__56_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__56_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__56_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__56_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__56_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__44_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__44_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__44_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__44_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__44_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__56_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__44_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_46_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__34_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__46_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__56_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__45_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__45_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__45_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__45_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__45_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__45_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__45_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__45_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__45_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__45_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__45_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__45_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__45_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__45_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__45_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__45_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__45_ccff_tail));

	tile_1__2_ tile_5__4_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__57_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__57_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__57_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__57_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__57_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__57_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__45_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__45_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__45_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__45_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__45_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__57_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__45_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_5__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__35_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__4_sb_1__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__35_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__46_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__46_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__46_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__46_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__46_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__46_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__46_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__46_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__46_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__46_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__46_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__46_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__46_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__46_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__46_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__46_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__46_ccff_tail));

	tile_1__2_ tile_5__7_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__58_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__58_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__58_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__58_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__58_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__58_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__58_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__6__4_cby_1__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_48_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__36_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__48_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[13]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__47_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__47_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__47_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__47_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__47_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__47_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__47_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__47_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__47_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__47_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__47_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__47_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__47_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__47_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__47_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__47_ccff_tail));

	tile_1__2_ tile_5__8_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__59_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__59_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__59_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__59_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__59_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__59_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__47_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__47_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__47_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__47_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__47_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__59_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__47_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_49_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__37_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__49_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[14]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__48_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__48_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__48_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__48_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__48_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__48_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__48_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__48_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__48_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__48_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__48_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__48_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__48_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__48_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__48_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__48_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__48_ccff_tail));

	tile_1__2_ tile_5__9_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__60_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__60_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__60_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__60_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__60_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__60_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__48_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__48_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__48_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__48_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__48_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__60_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__48_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_5__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__38_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__10__2_sb_1__9__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__60_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__49_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__49_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__49_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__49_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__49_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__49_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__49_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__49_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__49_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__49_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__49_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__49_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__49_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__49_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__49_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__49_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__49_ccff_tail));

	tile_1__2_ tile_5__12_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__61_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__61_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__61_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__61_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__61_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__61_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__61_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__11__2_cby_1__11__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_51_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__39_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__51_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__39_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__50_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__50_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__50_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__50_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__50_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__50_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__50_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__50_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__50_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__50_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__50_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__50_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__50_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__50_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__50_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__50_ccff_tail));

	tile_1__2_ tile_5__13_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__62_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__62_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__62_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__62_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__62_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__62_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__50_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__50_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__50_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__50_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__50_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__62_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__50_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_5__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__40_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__5_sb_1__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__62_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__51_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__51_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__51_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__51_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__51_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__51_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__51_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__51_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__51_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__51_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__51_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__51_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__51_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__51_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__51_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__51_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__51_ccff_tail));

	tile_1__2_ tile_5__16_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__63_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__63_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__63_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__63_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__63_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__63_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__63_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__6__5_cby_1__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_53_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__41_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__53_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__41_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__52_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__52_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__52_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__52_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__52_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__52_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__52_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__52_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__52_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__52_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__52_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__52_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__52_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__52_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__52_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[26]));

	tile_1__2_ tile_5__17_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__64_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__64_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__64_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__64_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__64_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__64_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__52_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__52_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__52_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__52_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__52_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__64_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__52_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_54_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__42_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__54_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__64_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__53_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__53_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__53_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__53_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__53_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__53_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__53_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__53_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__53_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__53_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__53_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__53_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__53_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__53_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__53_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__53_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__53_ccff_tail));

	tile_1__2_ tile_5__18_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__65_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__65_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__65_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__65_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__65_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__65_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__53_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__53_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__53_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__53_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__53_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__65_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__53_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__4_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_5__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__43_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__19__4_sb_1__18__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__43_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__54_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__54_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__54_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__54_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__54_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__54_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__54_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__54_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__54_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__54_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__54_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__54_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__54_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__54_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__54_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__54_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__54_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__54_ccff_tail));

	tile_1__2_ tile_6__2_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__66_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__66_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__66_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__66_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__66_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__66_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__66_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__1__5_cby_1__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_56_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__44_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__56_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[4]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__55_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__55_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__55_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__55_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__55_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__55_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__55_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__55_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__55_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__55_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__55_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__55_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__55_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__55_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__55_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__55_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__55_ccff_tail));

	tile_1__2_ tile_6__3_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__67_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__67_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__67_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__67_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__67_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__67_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__55_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__55_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__55_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__55_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__55_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__67_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__55_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_57_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__45_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__57_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__67_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__56_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__56_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__56_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__56_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__56_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__56_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__56_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__56_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__56_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__56_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__56_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__56_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__56_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__56_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__56_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__56_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__56_ccff_tail));

	tile_1__2_ tile_6__4_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__68_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__68_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__68_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__68_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__68_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__68_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__56_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__56_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__56_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__56_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__56_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__68_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__56_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_6__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__46_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__4_sb_2__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__46_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__57_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__57_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__57_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__57_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__57_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__57_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__57_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__57_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__57_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__57_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__57_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__57_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__57_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__57_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__57_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__57_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__57_ccff_tail));

	tile_1__2_ tile_6__7_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__69_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__69_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__69_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__69_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__69_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__69_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__69_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__6__4_cby_2__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_59_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__47_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__59_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__69_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__58_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__58_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__58_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__58_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__58_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__58_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__58_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__58_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__58_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__58_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__58_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__58_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__58_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__58_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__58_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[12]));

	tile_1__2_ tile_6__8_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__70_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__70_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__70_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__70_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__70_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__70_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__58_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__58_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__58_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__58_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__58_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__70_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__58_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_60_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__48_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__60_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__48_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__59_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__59_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__59_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__59_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__59_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__59_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__59_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__59_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__59_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__59_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__59_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__59_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__59_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__59_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__59_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__59_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__59_ccff_tail));

	tile_1__2_ tile_6__9_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__71_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__71_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__71_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__71_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__71_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__71_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__59_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__59_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__59_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__59_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__59_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__71_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__59_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_6__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__49_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__10__2_sb_2__9__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__71_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__60_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__60_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__60_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__60_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__60_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__60_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__60_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__60_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__60_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__60_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__60_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__60_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__60_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__60_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__60_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__60_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__60_ccff_tail));

	tile_1__2_ tile_6__12_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__72_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__72_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__72_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__72_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__72_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__72_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__72_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__11__2_cby_2__11__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_62_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__50_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__62_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__50_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__61_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__61_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__61_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__61_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__61_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__61_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__61_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__61_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__61_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__61_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__61_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__61_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__61_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__61_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__61_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__61_ccff_tail));

	tile_1__2_ tile_6__13_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__73_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__73_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__73_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__73_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__73_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__73_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__61_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__61_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__61_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__61_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__61_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__73_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__61_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_6__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__51_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__5_sb_2__4__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[23]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__62_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__62_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__62_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__62_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__62_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__62_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__62_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__62_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__62_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__62_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__62_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__62_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__62_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__62_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__62_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__62_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__62_ccff_tail));

	tile_1__2_ tile_6__16_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__74_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__74_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__74_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__74_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__74_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__74_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__74_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__6__5_cby_2__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_64_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__52_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__64_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[27]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__63_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__63_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__63_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__63_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__63_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__63_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__63_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__63_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__63_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__63_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__63_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__63_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__63_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__63_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__63_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__63_ccff_tail));

	tile_1__2_ tile_6__17_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__75_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__75_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__75_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__75_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__75_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__75_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__63_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__63_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__63_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__63_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__63_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__75_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__63_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_65_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__53_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__65_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__75_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__64_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__64_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__64_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__64_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__64_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__64_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__64_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__64_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__64_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__64_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__64_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__64_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__64_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__64_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__64_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__64_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__64_ccff_tail));

	tile_1__2_ tile_6__18_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__76_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__76_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__76_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__76_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__76_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__76_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__64_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__64_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__64_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__64_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__64_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__76_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__64_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__5_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_6__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__54_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__19__5_sb_1__18__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__54_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__65_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__65_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__65_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__65_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__65_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__65_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__65_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__65_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__65_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__65_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__65_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__65_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__65_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__65_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__65_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__65_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__65_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__65_ccff_tail));

	tile_1__2_ tile_7__2_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__77_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__77_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__77_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__77_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__77_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__77_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__77_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__1__6_cby_1__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_67_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__55_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__67_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__55_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__66_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__66_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__66_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__66_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__66_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__66_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__66_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__66_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__66_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__66_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__66_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__66_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__66_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__66_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__66_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__66_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__66_ccff_tail));

	tile_1__2_ tile_7__3_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__78_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__78_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__78_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__78_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__78_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__78_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__66_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__66_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__66_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__66_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__66_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__78_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__66_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_68_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__56_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__68_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__78_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__67_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__67_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__67_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__67_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__67_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__67_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__67_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__67_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__67_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__67_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__67_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__67_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__67_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__67_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__67_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__67_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__67_ccff_tail));

	tile_1__2_ tile_7__4_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__79_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__79_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__79_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__79_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__79_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__79_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__67_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__67_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__67_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__67_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__67_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__79_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__67_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_7__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__57_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__6_sb_1__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__57_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__68_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__68_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__68_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__68_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__68_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__68_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__68_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__68_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__68_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__68_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__68_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__68_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__68_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__68_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__68_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__68_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__68_ccff_tail));

	tile_1__2_ tile_7__7_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__80_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__80_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__80_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__80_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__80_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__80_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__80_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__6__6_cby_1__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_70_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__58_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__70_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__80_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__69_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__69_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__69_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__69_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__69_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__69_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__69_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__69_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__69_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__69_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__69_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__69_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__69_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__69_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__69_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__69_ccff_tail));

	tile_1__2_ tile_7__8_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__81_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__81_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__81_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__81_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__81_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__81_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__69_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__69_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__69_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__69_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__69_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__81_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__69_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_71_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__59_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__71_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__59_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__70_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__70_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__70_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__70_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__70_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__70_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__70_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__70_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__70_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__70_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__70_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__70_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__70_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__70_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__70_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__70_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__70_ccff_tail));

	tile_1__2_ tile_7__9_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__82_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__82_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__82_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__82_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__82_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__82_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__70_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__70_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__70_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__70_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__70_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__82_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__70_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_7__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__60_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__10__3_sb_1__9__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__82_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__71_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__71_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__71_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__71_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__71_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__71_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__71_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__71_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__71_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__71_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__71_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__71_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__71_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__71_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__71_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__71_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__71_ccff_tail));

	tile_1__2_ tile_7__12_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__83_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__83_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__83_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__83_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__83_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__83_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__83_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__11__3_cby_1__11__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_73_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__61_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__73_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__61_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__72_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__72_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__72_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__72_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__72_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__72_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__72_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__72_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__72_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__72_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__72_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__72_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__72_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__72_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__72_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__72_ccff_tail));

	tile_1__2_ tile_7__13_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__84_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__84_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__84_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__84_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__84_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__84_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__72_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__72_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__72_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__72_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__72_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__84_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__72_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_7__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__62_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__7_sb_1__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__84_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__73_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__73_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__73_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__73_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__73_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__73_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__73_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__73_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__73_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__73_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__73_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__73_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__73_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__73_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__73_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__73_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[22]));

	tile_1__2_ tile_7__16_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__85_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__85_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__85_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__85_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__85_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__85_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__85_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__6__7_cby_1__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_75_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__63_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__75_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__63_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__74_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__74_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__74_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__74_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__74_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__74_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__74_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__74_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__74_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__74_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__74_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__74_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__74_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__74_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__74_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__74_ccff_tail));

	tile_1__2_ tile_7__17_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__86_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__86_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__86_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__86_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__86_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__86_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__74_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__74_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__74_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__74_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__74_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__86_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__74_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_76_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__64_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__76_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__86_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__75_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__75_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__75_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__75_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__75_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__75_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__75_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__75_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__75_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__75_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__75_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__75_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__75_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__75_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__75_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__75_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__75_ccff_tail));

	tile_1__2_ tile_7__18_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__87_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__87_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__87_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__87_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__87_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__87_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__75_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__75_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__75_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__75_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__75_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__87_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__75_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__6_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_7__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__65_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__19__6_sb_1__18__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__65_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__76_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__76_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__76_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__76_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__76_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__76_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__76_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__76_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__76_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__76_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__76_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__76_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__76_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__76_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__76_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__76_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__76_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__76_ccff_tail));

	tile_1__2_ tile_8__2_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__88_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__88_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__88_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__88_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__88_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__88_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__88_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__1__7_cby_1__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_78_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__66_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__78_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__66_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__77_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__77_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__77_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__77_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__77_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__77_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__77_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__77_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__77_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__77_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__77_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__77_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__77_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__77_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__77_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__77_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__77_ccff_tail));

	tile_1__2_ tile_8__3_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__89_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__89_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__89_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__89_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__89_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__89_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__77_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__77_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__77_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__77_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__77_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__89_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__77_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_79_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__67_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__79_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__89_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__78_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__78_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__78_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__78_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__78_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__78_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__78_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__78_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__78_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__78_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__78_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__78_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__78_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__78_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__78_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__78_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__78_ccff_tail));

	tile_1__2_ tile_8__4_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__90_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__90_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__90_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__90_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__90_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__90_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__78_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__78_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__78_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__78_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__78_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__90_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__78_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_8__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__68_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__6_sb_2__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__68_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__79_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__79_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__79_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__79_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__79_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__79_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__79_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__79_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__79_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__79_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__79_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__79_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__79_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__79_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__79_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__79_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__79_ccff_tail));

	tile_1__2_ tile_8__7_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__91_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__91_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__91_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__91_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__91_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__91_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__91_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__6__6_cby_2__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_81_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__69_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__81_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__91_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__80_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__80_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__80_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__80_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__80_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__80_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__80_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__80_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__80_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__80_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__80_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__80_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__80_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__80_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__80_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__80_ccff_tail));

	tile_1__2_ tile_8__8_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__92_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__92_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__92_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__92_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__92_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__92_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__80_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__80_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__80_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__80_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__80_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__92_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__80_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_82_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__70_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__82_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__70_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__81_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__81_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__81_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__81_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__81_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__81_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__81_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__81_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__81_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__81_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__81_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__81_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__81_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__81_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__81_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__81_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__81_ccff_tail));

	tile_1__2_ tile_8__9_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__93_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__93_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__93_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__93_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__93_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__93_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__81_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__81_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__81_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__81_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__81_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__93_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__81_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_8__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__71_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__10__3_sb_2__9__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__93_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__82_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__82_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__82_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__82_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__82_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__82_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__82_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__82_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__82_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__82_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__82_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__82_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__82_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__82_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__82_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__82_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__82_ccff_tail));

	tile_1__2_ tile_8__12_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__94_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__94_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__94_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__94_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__94_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__94_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__94_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__11__3_cby_2__11__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_84_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__72_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__84_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__72_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__83_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__83_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__83_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__83_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__83_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__83_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__83_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__83_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__83_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__83_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__83_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__83_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__83_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__83_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__83_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__83_ccff_tail));

	tile_1__2_ tile_8__13_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__95_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__95_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__95_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__95_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__95_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__95_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__83_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__83_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__83_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__83_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__83_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__95_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__83_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_8__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__73_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__7_sb_2__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__95_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__84_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__84_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__84_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__84_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__84_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__84_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__84_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__84_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__84_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__84_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__84_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__84_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__84_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__84_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__84_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__84_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__84_ccff_tail));

	tile_1__2_ tile_8__16_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__96_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__96_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__96_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__96_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__96_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__96_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__96_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__6__7_cby_2__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_86_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__74_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__86_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__74_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__85_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__85_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__85_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__85_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__85_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__85_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__85_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__85_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__85_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__85_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__85_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__85_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__85_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__85_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__85_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__85_ccff_tail));

	tile_1__2_ tile_8__17_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__97_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__97_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__97_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__97_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__97_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__97_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__85_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__85_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__85_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__85_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__85_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__97_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__85_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_87_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__75_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__87_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__97_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__86_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__86_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__86_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__86_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__86_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__86_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__86_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__86_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__86_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__86_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__86_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__86_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__86_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__86_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__86_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__86_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__86_ccff_tail));

	tile_1__2_ tile_8__18_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__98_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__98_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__98_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__98_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__98_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__98_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__86_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__86_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__86_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__86_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__86_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__98_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__86_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__7_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_8__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__76_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__19__7_sb_1__18__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__76_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__87_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__87_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__87_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__87_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__87_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__87_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__87_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__87_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__87_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__87_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__87_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__87_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__87_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__87_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__87_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__87_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__87_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__87_ccff_tail));

	tile_1__2_ tile_9__2_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__99_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__99_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__99_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__99_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__99_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__99_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__99_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__1__8_cby_1__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_89_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__77_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__89_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__77_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__88_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__88_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__88_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__88_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__88_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__88_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__88_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__88_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__88_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__88_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__88_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__88_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__88_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__88_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__88_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__88_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__88_ccff_tail));

	tile_1__2_ tile_9__3_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__100_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__100_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__100_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__100_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__100_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__100_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__88_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__88_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__88_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__88_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__88_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__100_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__88_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_90_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__78_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__90_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__100_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__89_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__89_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__89_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__89_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__89_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__89_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__89_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__89_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__89_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__89_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__89_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__89_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__89_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__89_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__89_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__89_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__89_ccff_tail));

	tile_1__2_ tile_9__4_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__101_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__101_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__101_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__101_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__101_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__101_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__89_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__89_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__89_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__89_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__89_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__101_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__89_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_9__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__79_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__8_sb_1__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__79_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__90_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__90_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__90_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__90_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__90_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__90_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__90_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__90_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__90_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__90_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__90_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__90_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__90_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__90_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__90_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__90_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[7]));

	tile_1__2_ tile_9__7_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__102_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__102_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__102_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__102_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__102_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__102_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__102_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__6__8_cby_1__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_92_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__80_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__92_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__102_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__91_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__91_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__91_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__91_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__91_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__91_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__91_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__91_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__91_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__91_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__91_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__91_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__91_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__91_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__91_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__91_ccff_tail));

	tile_1__2_ tile_9__8_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__103_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__103_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__103_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__103_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__103_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__103_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__91_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__91_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__91_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__91_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__91_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__103_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__91_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_93_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__81_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__93_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__81_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__92_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__92_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__92_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__92_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__92_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__92_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__92_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__92_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__92_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__92_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__92_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__92_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__92_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__92_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__92_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__92_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__92_ccff_tail));

	tile_1__2_ tile_9__9_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__104_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__104_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__104_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__104_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__104_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__104_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__92_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__92_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__92_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__92_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__92_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__104_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__92_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_9__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__82_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__10__4_sb_1__9__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__104_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__93_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__93_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__93_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__93_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__93_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__93_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__93_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__93_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__93_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__93_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__93_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__93_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__93_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__93_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__93_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__93_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__93_ccff_tail));

	tile_1__2_ tile_9__12_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__105_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__105_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__105_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__105_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__105_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__105_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__105_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__11__4_cby_1__11__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_95_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__83_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__95_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__83_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__94_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__94_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__94_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__94_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__94_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__94_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__94_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__94_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__94_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__94_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__94_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__94_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__94_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__94_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__94_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__94_ccff_tail));

	tile_1__2_ tile_9__13_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__106_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__106_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__106_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__106_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__106_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__106_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__94_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__94_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__94_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__94_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__94_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__106_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__94_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_9__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__84_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__9_sb_1__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__106_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__95_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__95_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__95_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__95_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__95_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__95_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__95_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__95_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__95_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__95_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__95_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__95_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__95_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__95_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__95_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__95_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__95_ccff_tail));

	tile_1__2_ tile_9__16_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__107_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__107_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__107_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__107_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__107_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__107_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__107_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__6__9_cby_1__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_97_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__85_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__97_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__85_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__96_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__96_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__96_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__96_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__96_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__96_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__96_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__96_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__96_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__96_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__96_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__96_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__96_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__96_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__96_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__96_ccff_tail));

	tile_1__2_ tile_9__17_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__108_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__108_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__108_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__108_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__108_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__108_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__96_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__96_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__96_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__96_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__96_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__108_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__96_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_98_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__86_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__98_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__108_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__97_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__97_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__97_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__97_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__97_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__97_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__97_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__97_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__97_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__97_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__97_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__97_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__97_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__97_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__97_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__97_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__97_ccff_tail));

	tile_1__2_ tile_9__18_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__109_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__109_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__109_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__109_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__109_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__109_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__97_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__97_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__97_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__97_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__97_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__109_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__97_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__8_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_9__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__87_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__19__8_sb_1__18__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__87_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__98_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__98_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__98_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__98_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__98_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__98_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__98_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__98_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__98_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__98_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__98_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__98_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__98_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__98_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__98_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__98_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__98_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[30]));

	tile_1__2_ tile_10__2_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__110_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__110_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__110_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__110_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__110_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__110_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__110_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__1__9_cby_1__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_100_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__88_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__100_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__88_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__99_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__99_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__99_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__99_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__99_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__99_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__99_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__99_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__99_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__99_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__99_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__99_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__99_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__99_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__99_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__99_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__99_ccff_tail));

	tile_1__2_ tile_10__3_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__111_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__111_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__111_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__111_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__111_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__111_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__99_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__99_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__99_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__99_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__99_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__111_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__99_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_101_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__89_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__101_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__111_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__100_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__100_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__100_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__100_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__100_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__100_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__100_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__100_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__100_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__100_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__100_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__100_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__100_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__100_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__100_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__100_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__100_ccff_tail));

	tile_1__2_ tile_10__4_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__112_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__112_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__112_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__112_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__112_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__112_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__100_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__100_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__100_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__100_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__100_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__112_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__100_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_10__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__90_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__8_sb_2__4__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[8]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__101_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__101_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__101_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__101_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__101_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__101_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__101_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__101_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__101_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__101_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__101_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__101_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__101_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__101_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__101_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__101_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__101_ccff_tail));

	tile_1__2_ tile_10__7_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__113_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__113_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__113_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__113_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__113_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__113_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__113_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__6__8_cby_2__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_103_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__91_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__103_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__113_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__102_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__102_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__102_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__102_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__102_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__102_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__102_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__102_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__102_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__102_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__102_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__102_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__102_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__102_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__102_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__102_ccff_tail));

	tile_1__2_ tile_10__8_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__114_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__114_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__114_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__114_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__114_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__114_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__102_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__102_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__102_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__102_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__102_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__114_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__102_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_104_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__92_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__104_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__92_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__103_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__103_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__103_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__103_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__103_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__103_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__103_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__103_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__103_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__103_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__103_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__103_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__103_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__103_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__103_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__103_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__103_ccff_tail));

	tile_1__2_ tile_10__9_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__115_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__115_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__115_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__115_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__115_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__115_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__103_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__103_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__103_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__103_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__103_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__115_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__103_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_10__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__93_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__10__4_sb_2__9__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__115_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__104_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__104_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__104_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__104_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__104_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__104_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__104_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__104_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__104_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__104_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__104_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__104_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__104_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__104_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__104_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__104_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__104_ccff_tail));

	tile_1__2_ tile_10__12_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__116_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__116_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__116_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__116_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__116_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__116_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__116_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__11__4_cby_2__11__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_106_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__94_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__106_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__94_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__105_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__105_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__105_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__105_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__105_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__105_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__105_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__105_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__105_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__105_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__105_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__105_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__105_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__105_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__105_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[20]));

	tile_1__2_ tile_10__13_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__117_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__117_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__117_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__117_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__117_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__117_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__105_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__105_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__105_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__105_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__105_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__117_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__105_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_10__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__95_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__9_sb_2__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__117_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__106_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__106_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__106_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__106_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__106_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__106_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__106_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__106_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__106_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__106_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__106_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__106_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__106_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__106_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__106_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__106_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__106_ccff_tail));

	tile_1__2_ tile_10__16_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__118_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__118_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__118_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__118_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__118_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__118_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__118_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__6__9_cby_2__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_108_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__96_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__108_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__96_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__107_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__107_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__107_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__107_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__107_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__107_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__107_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__107_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__107_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__107_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__107_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__107_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__107_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__107_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__107_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__107_ccff_tail));

	tile_1__2_ tile_10__17_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__119_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__119_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__119_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__119_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__119_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__119_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__107_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__107_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__107_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__107_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__107_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__119_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__107_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_109_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__97_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__109_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__119_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__108_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__108_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__108_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__108_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__108_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__108_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__108_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__108_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__108_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__108_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__108_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__108_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__108_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__108_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__108_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__108_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__108_ccff_tail));

	tile_1__2_ tile_10__18_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__120_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__120_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__120_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__120_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__120_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__120_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__108_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__108_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__108_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__108_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__108_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__120_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__108_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__9_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_10__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__98_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__19__9_sb_1__18__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[31]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__109_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__109_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__109_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__109_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__109_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__109_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__109_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__109_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__109_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__109_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__109_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__109_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__109_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__109_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__109_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__109_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__109_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__109_ccff_tail));

	tile_1__2_ tile_11__2_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__121_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__121_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__121_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__121_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__121_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__121_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__121_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__1__10_cby_1__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_111_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__99_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__111_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__99_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__110_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__110_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__110_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__110_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__110_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__110_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__110_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__110_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__110_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__110_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__110_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__110_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__110_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__110_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__110_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__110_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__110_ccff_tail));

	tile_1__2_ tile_11__3_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__122_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__122_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__122_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__122_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__122_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__122_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__110_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__110_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__110_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__110_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__110_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__122_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__110_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_112_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__100_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__112_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[6]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__111_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__111_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__111_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__111_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__111_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__111_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__111_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__111_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__111_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__111_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__111_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__111_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__111_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__111_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__111_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__111_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__111_ccff_tail));

	tile_1__2_ tile_11__4_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__123_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__123_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__123_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__123_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__123_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__123_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__111_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__111_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__111_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__111_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__111_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__123_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__111_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_11__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__101_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__10_sb_1__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__101_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__112_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__112_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__112_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__112_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__112_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__112_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__112_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__112_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__112_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__112_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__112_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__112_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__112_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__112_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__112_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__112_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__112_ccff_tail));

	tile_1__2_ tile_11__7_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__124_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__124_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__124_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__124_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__124_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__124_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__124_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__6__10_cby_1__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_114_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__102_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__114_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__124_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__113_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__113_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__113_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__113_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__113_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__113_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__113_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__113_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__113_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__113_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__113_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__113_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__113_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__113_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__113_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__113_ccff_tail));

	tile_1__2_ tile_11__8_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__125_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__125_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__125_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__125_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__125_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__125_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__113_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__113_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__113_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__113_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__113_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__125_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__113_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_115_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__103_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__115_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__103_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__114_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__114_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__114_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__114_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__114_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__114_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__114_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__114_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__114_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__114_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__114_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__114_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__114_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__114_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__114_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__114_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__114_ccff_tail));

	tile_1__2_ tile_11__9_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__126_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__126_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__126_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__126_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__126_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__126_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__114_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__114_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__114_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__114_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__114_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__126_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__114_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_11__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__104_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__10__5_sb_1__9__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__126_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__115_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__115_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__115_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__115_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__115_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__115_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__115_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__115_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__115_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__115_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__115_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__115_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__115_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__115_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__115_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__115_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__115_ccff_tail));

	tile_1__2_ tile_11__12_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__127_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__127_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__127_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__127_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__127_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__127_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__127_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__11__5_cby_1__11__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_117_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__105_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__117_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[21]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__116_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__116_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__116_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__116_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__116_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__116_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__116_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__116_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__116_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__116_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__116_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__116_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__116_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__116_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__116_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__116_ccff_tail));

	tile_1__2_ tile_11__13_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__128_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__128_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__128_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__128_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__128_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__128_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__116_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__116_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__116_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__116_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__116_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__128_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__116_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_11__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__106_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__11_sb_1__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__128_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__117_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__117_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__117_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__117_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__117_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__117_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__117_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__117_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__117_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__117_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__117_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__117_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__117_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__117_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__117_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__117_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__117_ccff_tail));

	tile_1__2_ tile_11__16_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__129_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__129_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__129_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__129_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__129_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__129_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__129_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__6__11_cby_1__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_119_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__107_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__119_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__107_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__118_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__118_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__118_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__118_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__118_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__118_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__118_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__118_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__118_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__118_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__118_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__118_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__118_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__118_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__118_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__118_ccff_tail));

	tile_1__2_ tile_11__17_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__130_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__130_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__130_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__130_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__130_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__130_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__118_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__118_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__118_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__118_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__118_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__130_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__118_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_120_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__108_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__120_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[29]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__119_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__119_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__119_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__119_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__119_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__119_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__119_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__119_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__119_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__119_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__119_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__119_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__119_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__119_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__119_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__119_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__119_ccff_tail));

	tile_1__2_ tile_11__18_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__131_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__131_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__131_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__131_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__131_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__131_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__119_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__119_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__119_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__119_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__119_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__131_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__119_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__10_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_11__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__109_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__19__10_sb_1__18__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__109_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__120_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__120_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__120_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__120_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__120_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__120_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__120_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__120_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__120_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__120_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__120_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__120_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__120_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__120_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__120_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__120_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__120_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__120_ccff_tail));

	tile_1__2_ tile_12__2_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__132_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__132_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__132_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__132_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__132_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__132_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__132_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__1__11_cby_1__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_122_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__110_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__122_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__110_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__121_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__121_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__121_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__121_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__121_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__121_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__121_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__121_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__121_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__121_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__121_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__121_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__121_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__121_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__121_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__121_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__121_ccff_tail));

	tile_1__2_ tile_12__3_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__133_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__133_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__133_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__133_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__133_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__133_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__121_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__121_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__121_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__121_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__121_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__133_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__121_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_123_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__111_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__123_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__133_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__122_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__122_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__122_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__122_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__122_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__122_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__122_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__122_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__122_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__122_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__122_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__122_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__122_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__122_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__122_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__122_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[5]));

	tile_1__2_ tile_12__4_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__134_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__134_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__134_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__134_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__134_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__134_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__122_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__122_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__122_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__122_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__122_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__134_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__122_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_12__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__112_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__10_sb_2__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__112_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__123_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__123_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__123_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__123_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__123_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__123_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__123_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__123_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__123_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__123_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__123_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__123_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__123_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__123_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__123_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__123_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__123_ccff_tail));

	tile_1__2_ tile_12__7_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__135_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__135_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__135_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__135_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__135_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__135_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__135_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__6__10_cby_2__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_125_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__113_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__125_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__135_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__124_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__124_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__124_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__124_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__124_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__124_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__124_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__124_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__124_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__124_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__124_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__124_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__124_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__124_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__124_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__124_ccff_tail));

	tile_1__2_ tile_12__8_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__136_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__136_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__136_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__136_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__136_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__136_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__124_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__124_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__124_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__124_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__124_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__136_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__124_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_126_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__114_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__126_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__114_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__125_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__125_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__125_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__125_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__125_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__125_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__125_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__125_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__125_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__125_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__125_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__125_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__125_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__125_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__125_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__125_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__125_ccff_tail));

	tile_1__2_ tile_12__9_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__137_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__137_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__137_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__137_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__137_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__137_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__125_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__125_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__125_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__125_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__125_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__137_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__125_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_12__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__115_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__10__5_sb_2__9__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[16]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__126_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__126_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__126_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__126_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__126_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__126_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__126_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__126_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__126_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__126_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__126_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__126_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__126_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__126_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__126_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__126_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__126_ccff_tail));

	tile_1__2_ tile_12__12_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__138_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__138_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__138_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__138_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__138_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__138_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__138_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__11__5_cby_2__11__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_128_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__116_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__128_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__116_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__127_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__127_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__127_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__127_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__127_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__127_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__127_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__127_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__127_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__127_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__127_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__127_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__127_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__127_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__127_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__127_ccff_tail));

	tile_1__2_ tile_12__13_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__139_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__139_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__139_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__139_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__139_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__139_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__127_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__127_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__127_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__127_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__127_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__139_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__127_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_12__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__117_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__11_sb_2__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__139_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__128_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__128_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__128_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__128_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__128_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__128_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__128_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__128_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__128_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__128_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__128_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__128_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__128_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__128_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__128_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__128_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__128_ccff_tail));

	tile_1__2_ tile_12__16_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__140_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__140_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__140_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__140_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__140_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__140_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__140_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__6__11_cby_2__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_130_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__118_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__130_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__118_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__129_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__129_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__129_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__129_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__129_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__129_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__129_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__129_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__129_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__129_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__129_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__129_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__129_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__129_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__129_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__129_ccff_tail));

	tile_1__2_ tile_12__17_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__141_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__141_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__141_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__141_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__141_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__141_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__129_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__129_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__129_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__129_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__129_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__141_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__129_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_131_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__119_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__131_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__141_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__130_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__130_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__130_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__130_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__130_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__130_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__130_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__130_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__130_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__130_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__130_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__130_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__130_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__130_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__130_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__130_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[28]));

	tile_1__2_ tile_12__18_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__142_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__142_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__142_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__142_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__142_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__142_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__130_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__130_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__130_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__130_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__130_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__142_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__130_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__11_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_12__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__120_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__19__11_sb_1__18__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__120_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__131_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__131_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__131_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__131_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__131_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__131_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__131_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__131_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__131_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__131_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__131_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__131_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__131_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__131_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__131_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__131_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__131_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__131_ccff_tail));

	tile_1__2_ tile_13__2_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__143_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__143_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__143_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__143_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__143_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__143_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__143_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__1__12_cby_1__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_133_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__121_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__133_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__121_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__132_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__132_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__132_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__132_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__132_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__132_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__132_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__132_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__132_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__132_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__132_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__132_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__132_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__132_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__132_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__132_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__132_ccff_tail));

	tile_1__2_ tile_13__3_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__144_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__144_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__144_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__144_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__144_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__144_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__132_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__132_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__132_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__132_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__132_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__144_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__132_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_134_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__122_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__134_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__144_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__133_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__133_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__133_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__133_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__133_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__133_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__133_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__133_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__133_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__133_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__133_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__133_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__133_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__133_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__133_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__133_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__133_ccff_tail));

	tile_1__2_ tile_13__4_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__145_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__145_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__145_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__145_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__145_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__145_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__133_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__133_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__133_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__133_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__133_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__145_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__133_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_13__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__123_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__12_sb_1__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__123_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__134_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__134_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__134_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__134_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__134_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__134_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__134_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__134_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__134_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__134_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__134_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__134_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__134_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__134_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__134_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__134_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__134_ccff_tail));

	tile_1__2_ tile_13__7_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__146_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__146_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__146_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__146_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__146_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__146_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__146_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__6__12_cby_1__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_136_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__124_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__136_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__146_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__135_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__135_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__135_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__135_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__135_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__135_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__135_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__135_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__135_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__135_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__135_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__135_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__135_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__135_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__135_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__135_ccff_tail));

	tile_1__2_ tile_13__8_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__147_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__147_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__147_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__147_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__147_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__147_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__135_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__135_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__135_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__135_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__135_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__147_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__135_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_137_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__125_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__137_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__125_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__136_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__136_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__136_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__136_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__136_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__136_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__136_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__136_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__136_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__136_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__136_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__136_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__136_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__136_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__136_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__136_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__136_ccff_tail));

	tile_1__2_ tile_13__9_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__148_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__148_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__148_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__148_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__148_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__148_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__136_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__136_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__136_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__136_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__136_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__148_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__136_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_13__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__126_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__10__6_sb_1__9__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__148_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__137_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__137_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__137_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__137_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__137_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__137_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__137_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__137_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__137_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__137_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__137_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__137_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__137_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__137_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__137_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__137_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[15]));

	tile_1__2_ tile_13__12_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__149_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__149_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__149_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__149_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__149_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__149_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__149_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__11__6_cby_1__11__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_139_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__127_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__139_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__127_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__138_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__138_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__138_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__138_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__138_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__138_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__138_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__138_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__138_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__138_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__138_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__138_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__138_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__138_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__138_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__138_ccff_tail));

	tile_1__2_ tile_13__13_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__150_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__150_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__150_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__150_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__150_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__150_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__138_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__138_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__138_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__138_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__138_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__150_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__138_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_13__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__128_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__13_sb_1__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__150_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__139_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__139_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__139_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__139_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__139_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__139_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__139_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__139_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__139_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__139_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__139_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__139_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__139_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__139_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__139_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__139_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__139_ccff_tail));

	tile_1__2_ tile_13__16_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__151_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__151_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__151_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__151_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__151_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__151_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__151_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__6__13_cby_1__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_141_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__129_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__141_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__129_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__140_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__140_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__140_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__140_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__140_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__140_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__140_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__140_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__140_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__140_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__140_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__140_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__140_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__140_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__140_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__140_ccff_tail));

	tile_1__2_ tile_13__17_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__152_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__152_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__152_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__152_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__152_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__152_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__140_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__140_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__140_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__140_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__140_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__152_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__140_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_142_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__130_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__142_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__152_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__141_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__141_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__141_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__141_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__141_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__141_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__141_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__141_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__141_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__141_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__141_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__141_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__141_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__141_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__141_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__141_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__141_ccff_tail));

	tile_1__2_ tile_13__18_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__153_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__153_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__153_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__153_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__153_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__153_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__141_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__141_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__141_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__141_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__141_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__153_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__141_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__12_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_13__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__131_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__19__12_sb_1__18__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__131_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__142_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__142_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__142_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__142_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__142_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__142_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__142_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__142_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__142_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__142_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__142_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__142_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__142_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__142_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__142_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__142_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__142_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__142_ccff_tail));

	tile_1__2_ tile_14__2_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__154_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__154_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__154_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__154_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__154_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__154_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__154_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__1__13_cby_1__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_144_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__132_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__144_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__132_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__143_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__143_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__143_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__143_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__143_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__143_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__143_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__143_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__143_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__143_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__143_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__143_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__143_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__143_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__143_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__143_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__143_ccff_tail));

	tile_1__2_ tile_14__3_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__155_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__155_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__155_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__155_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__155_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__155_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__143_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__143_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__143_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__143_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__143_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__155_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__143_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_145_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__133_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__145_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__155_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__144_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__144_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__144_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__144_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__144_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__144_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__144_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__144_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__144_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__144_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__144_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__144_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__144_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__144_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__144_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__144_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__144_ccff_tail));

	tile_1__2_ tile_14__4_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__156_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__156_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__156_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__156_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__156_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__156_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__144_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__144_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__144_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__144_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__144_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__156_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__144_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_14__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__134_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__12_sb_2__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__134_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__145_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__145_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__145_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__145_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__145_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__145_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__145_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__145_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__145_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__145_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__145_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__145_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__145_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__145_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__145_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__145_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__145_ccff_tail));

	tile_1__2_ tile_14__7_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__157_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__157_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__157_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__157_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__157_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__157_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__157_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__6__12_cby_2__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_147_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__135_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__147_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__157_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__146_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__146_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__146_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__146_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__146_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__146_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__146_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__146_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__146_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__146_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__146_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__146_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__146_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__146_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__146_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__146_ccff_tail));

	tile_1__2_ tile_14__8_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__158_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__158_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__158_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__158_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__158_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__158_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__146_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__146_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__146_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__146_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__146_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__158_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__146_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_148_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__136_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__148_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__136_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__147_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__147_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__147_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__147_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__147_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__147_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__147_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__147_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__147_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__147_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__147_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__147_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__147_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__147_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__147_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__147_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__147_ccff_tail));

	tile_1__2_ tile_14__9_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__159_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__159_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__159_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__159_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__159_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__159_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__147_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__147_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__147_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__147_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__147_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__159_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__147_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_14__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__137_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__10__6_sb_2__9__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__159_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__148_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__148_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__148_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__148_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__148_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__148_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__148_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__148_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__148_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__148_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__148_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__148_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__148_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__148_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__148_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__148_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__148_ccff_tail));

	tile_1__2_ tile_14__12_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__160_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__160_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__160_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__160_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__160_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__160_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__160_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__11__6_cby_2__11__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_150_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__138_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__150_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__138_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__149_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__149_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__149_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__149_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__149_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__149_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__149_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__149_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__149_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__149_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__149_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__149_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__149_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__149_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__149_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__149_ccff_tail));

	tile_1__2_ tile_14__13_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__161_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__161_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__161_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__161_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__161_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__161_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__149_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__149_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__149_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__149_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__149_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__161_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__149_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_14__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__139_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__13_sb_2__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__161_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__150_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__150_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__150_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__150_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__150_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__150_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__150_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__150_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__150_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__150_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__150_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__150_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__150_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__150_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__150_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__150_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__150_ccff_tail));

	tile_1__2_ tile_14__16_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__162_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__162_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__162_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__162_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__162_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__162_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__162_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__6__13_cby_2__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_152_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__140_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__152_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__140_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__151_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__151_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__151_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__151_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__151_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__151_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__151_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__151_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__151_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__151_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__151_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__151_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__151_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__151_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__151_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__151_ccff_tail));

	tile_1__2_ tile_14__17_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__163_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__163_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__163_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__163_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__163_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__163_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__151_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__151_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__151_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__151_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__151_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__163_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__151_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_153_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__141_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__153_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__163_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__152_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__152_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__152_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__152_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__152_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__152_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__152_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__152_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__152_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__152_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__152_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__152_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__152_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__152_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__152_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__152_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__152_ccff_tail));

	tile_1__2_ tile_14__18_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__164_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__164_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__164_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__164_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__164_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__164_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__152_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__152_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__152_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__152_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__152_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__164_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__152_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__13_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_14__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__142_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__19__13_sb_1__18__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__142_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__153_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__153_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__153_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__153_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__153_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__153_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__153_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__153_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__153_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__153_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__153_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__153_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__153_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__153_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__153_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__153_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__153_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__153_ccff_tail));

	tile_1__2_ tile_15__2_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__165_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__165_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__165_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__165_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__165_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__165_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__165_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__1__14_cby_1__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_155_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__143_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__155_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__143_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__154_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__154_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__154_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__154_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__154_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__154_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__154_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__154_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__154_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__154_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__154_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__154_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__154_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__154_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__154_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__154_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__154_ccff_tail));

	tile_1__2_ tile_15__3_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__166_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__166_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__166_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__166_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__166_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__166_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__154_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__154_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__154_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__154_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__154_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__166_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__154_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_156_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__144_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__156_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__166_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__155_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__155_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__155_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__155_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__155_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__155_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__155_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__155_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__155_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__155_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__155_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__155_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__155_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__155_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__155_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__155_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__155_ccff_tail));

	tile_1__2_ tile_15__4_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__167_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__167_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__167_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__167_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__167_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__167_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__155_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__155_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__155_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__155_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__155_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__167_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__155_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_15__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__145_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__14_sb_1__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__145_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__156_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__156_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__156_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__156_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__156_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__156_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__156_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__156_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__156_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__156_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__156_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__156_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__156_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__156_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__156_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__156_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__156_ccff_tail));

	tile_1__2_ tile_15__7_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__168_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__168_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__168_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__168_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__168_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__168_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__168_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__6__14_cby_1__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_158_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__146_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__158_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__168_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__157_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__157_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__157_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__157_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__157_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__157_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__157_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__157_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__157_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__157_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__157_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__157_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__157_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__157_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__157_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__157_ccff_tail));

	tile_1__2_ tile_15__8_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__169_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__169_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__169_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__169_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__169_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__169_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__157_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__157_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__157_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__157_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__157_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__169_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__157_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_159_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__147_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__159_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__147_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__158_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__158_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__158_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__158_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__158_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__158_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__158_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__158_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__158_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__158_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__158_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__158_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__158_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__158_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__158_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__158_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[14]));

	tile_1__2_ tile_15__9_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__170_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__170_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__170_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__170_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__170_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__170_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__158_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__158_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__158_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__158_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__158_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__170_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__158_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_15__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__148_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__10__7_sb_1__9__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__170_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__159_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__159_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__159_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__159_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__159_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__159_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__159_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__159_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__159_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__159_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__159_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__159_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__159_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__159_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__159_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__159_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__159_ccff_tail));

	tile_1__2_ tile_15__12_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__171_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__171_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__171_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__171_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__171_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__171_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__171_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__11__7_cby_1__11__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_161_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__149_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__161_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__149_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__160_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__160_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__160_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__160_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__160_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__160_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__160_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__160_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__160_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__160_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__160_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__160_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__160_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__160_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__160_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__160_ccff_tail));

	tile_1__2_ tile_15__13_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__172_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__172_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__172_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__172_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__172_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__172_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__160_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__160_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__160_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__160_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__160_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__172_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__160_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_15__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__150_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__15_sb_1__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__172_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__161_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__161_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__161_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__161_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__161_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__161_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__161_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__161_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__161_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__161_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__161_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__161_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__161_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__161_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__161_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__161_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__161_ccff_tail));

	tile_1__2_ tile_15__16_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__173_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__173_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__173_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__173_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__173_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__173_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__173_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__6__15_cby_1__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_163_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__151_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__163_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__151_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__162_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__162_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__162_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__162_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__162_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__162_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__162_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__162_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__162_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__162_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__162_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__162_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__162_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__162_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__162_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__162_ccff_tail));

	tile_1__2_ tile_15__17_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__174_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__174_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__174_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__174_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__174_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__174_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__162_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__162_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__162_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__162_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__162_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__174_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__162_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_164_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__152_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__164_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__174_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__163_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__163_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__163_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__163_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__163_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__163_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__163_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__163_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__163_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__163_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__163_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__163_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__163_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__163_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__163_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__163_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__163_ccff_tail));

	tile_1__2_ tile_15__18_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__175_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__175_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__175_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__175_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__175_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__175_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__163_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__163_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__163_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__163_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__163_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__175_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__163_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__14_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_15__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__153_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__19__14_sb_1__18__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__153_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__164_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__164_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__164_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__164_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__164_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__164_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__164_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__164_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__164_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__164_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__164_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__164_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__164_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__164_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__164_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__164_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__164_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__164_ccff_tail));

	tile_1__2_ tile_16__2_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__176_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__176_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__176_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__176_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__176_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__176_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__176_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__1__15_cby_1__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_166_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__154_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__166_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__154_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__165_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__165_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__165_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__165_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__165_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__165_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__165_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__165_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__165_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__165_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__165_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__165_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__165_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__165_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__165_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__165_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[4]));

	tile_1__2_ tile_16__3_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__177_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__177_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__177_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__177_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__177_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__177_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__165_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__165_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__165_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__165_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__165_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__177_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__165_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_167_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__155_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__167_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__177_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__166_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__166_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__166_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__166_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__166_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__166_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__166_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__166_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__166_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__166_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__166_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__166_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__166_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__166_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__166_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__166_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__166_ccff_tail));

	tile_1__2_ tile_16__4_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__178_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__178_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__178_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__178_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__178_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__178_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__166_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__166_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__166_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__166_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__166_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__178_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__166_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_16__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__156_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__14_sb_2__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__156_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__167_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__167_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__167_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__167_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__167_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__167_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__167_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__167_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__167_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__167_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__167_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__167_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__167_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__167_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__167_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__167_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__167_ccff_tail));

	tile_1__2_ tile_16__7_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__179_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__179_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__179_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__179_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__179_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__179_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__179_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__6__14_cby_2__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_169_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__157_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__169_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[12]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__168_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__168_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__168_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__168_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__168_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__168_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__168_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__168_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__168_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__168_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__168_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__168_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__168_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__168_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__168_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__168_ccff_tail));

	tile_1__2_ tile_16__8_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__180_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__180_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__180_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__180_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__180_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__180_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__168_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__168_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__168_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__168_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__168_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__180_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__168_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_170_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__158_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__170_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[15]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__169_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__169_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__169_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__169_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__169_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__169_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__169_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__169_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__169_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__169_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__169_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__169_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__169_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__169_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__169_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__169_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__169_ccff_tail));

	tile_1__2_ tile_16__9_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__181_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__181_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__181_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__181_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__181_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__181_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__169_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__169_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__169_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__169_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__169_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__181_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__169_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_16__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__159_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__10__7_sb_2__9__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__181_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__170_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__170_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__170_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__170_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__170_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__170_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__170_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__170_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__170_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__170_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__170_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__170_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__170_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__170_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__170_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__170_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__170_ccff_tail));

	tile_1__2_ tile_16__12_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__182_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__182_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__182_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__182_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__182_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__182_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__182_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__11__7_cby_2__11__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_172_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__160_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__172_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__160_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__171_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__171_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__171_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__171_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__171_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__171_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__171_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__171_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__171_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__171_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__171_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__171_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__171_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__171_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__171_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__171_ccff_tail));

	tile_1__2_ tile_16__13_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__183_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__183_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__183_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__183_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__183_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__183_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__171_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__171_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__171_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__171_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__171_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__183_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__171_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_16__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__161_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__5__15_sb_2__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__183_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__172_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__172_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__172_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__172_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__172_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__172_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__172_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__172_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__172_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__172_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__172_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__172_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__172_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__172_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__172_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__172_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__172_ccff_tail));

	tile_1__2_ tile_16__16_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__184_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__184_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__184_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__184_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__184_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__184_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__184_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_2__6__15_cby_2__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_174_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__162_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__174_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__162_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__173_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__173_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__173_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__173_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__173_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__173_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__173_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__173_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__173_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__173_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__173_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__173_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__173_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__173_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__173_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[27]));

	tile_1__2_ tile_16__17_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__185_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__185_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__185_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__185_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__185_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__185_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__173_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__173_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__173_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__173_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__173_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__185_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__173_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_175_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__163_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__175_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__185_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__174_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__174_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__174_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__174_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__174_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__174_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__174_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__174_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__174_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__174_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__174_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__174_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__174_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__174_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__174_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__174_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__174_ccff_tail));

	tile_1__2_ tile_16__18_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__186_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__186_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__186_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__186_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__186_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__186_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__174_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__174_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__174_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__174_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__174_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_1__2__186_cbx_1__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__174_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__15_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_16__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__164_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__19__15_sb_1__18__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__164_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__175_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__175_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__175_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__175_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__175_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__175_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__175_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__175_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__175_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__175_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__175_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__175_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__175_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__175_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__175_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__175_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__175_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__175_ccff_tail));

	tile_1__2_ tile_17__2_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_18__2__0_cbx_18__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__1__16_cby_1__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_177_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__165_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__177_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[5]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__176_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__176_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__176_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__176_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__176_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__176_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__176_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__176_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__176_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__176_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__176_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__176_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__176_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__176_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__176_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__176_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__176_ccff_tail));

	tile_1__2_ tile_17__3_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__176_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__176_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__176_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__176_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__176_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_18__2__1_cbx_18__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__176_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_178_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__166_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__178_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_18__2__1_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__177_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__177_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__177_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__177_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__177_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__177_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__177_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__177_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__177_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__177_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__177_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__177_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__177_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__177_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__177_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__177_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__177_ccff_tail));

	tile_1__2_ tile_17__4_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__177_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__177_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__177_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__177_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__177_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_18__2__2_cbx_18__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__177_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_17__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__167_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_17__5__0_sb_17__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__167_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__178_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__178_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__178_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__178_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__178_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__178_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__178_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__178_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__178_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__178_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__178_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__178_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__178_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__178_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__178_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__178_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__178_ccff_tail));

	tile_1__2_ tile_17__7_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_18__2__3_cbx_18__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__6__16_cby_1__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_180_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__168_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__180_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_18__2__3_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__179_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__179_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__179_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__179_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__179_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__179_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__179_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__179_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__179_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__179_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__179_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__179_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__179_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__179_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__179_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[11]));

	tile_1__2_ tile_17__8_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__179_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__179_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__179_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__179_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__179_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_18__2__4_cbx_18__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__179_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_181_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__169_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__181_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__169_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__180_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__180_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__180_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__180_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__180_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__180_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__180_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__180_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__180_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__180_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__180_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__180_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__180_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__180_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__180_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__180_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__180_ccff_tail));

	tile_1__2_ tile_17__9_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__180_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__180_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__180_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__180_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__180_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_18__2__5_cbx_18__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__180_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_17__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__170_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_17__10__0_sb_17__9__chany_bottom_out[0:64]),
		.ccff_head(tile_18__2__5_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__181_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__181_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__181_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__181_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__181_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__181_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__181_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__181_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__181_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__181_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__181_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__181_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__181_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__181_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__181_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__181_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__181_ccff_tail));

	tile_1__2_ tile_17__12_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__11__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__11__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__11__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__11__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_18__2__6_cbx_18__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__11__8_cby_1__11__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_183_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__171_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__183_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__171_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__182_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__182_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__182_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__182_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__182_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__182_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__182_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__182_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__182_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__182_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__182_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__182_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__182_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__182_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__182_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__182_ccff_tail));

	tile_1__2_ tile_17__13_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__182_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__182_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__182_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__182_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__182_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_18__2__7_cbx_18__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__182_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_17__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__172_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_17__5__1_sb_17__4__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[22]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__183_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__183_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__183_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__183_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__183_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__183_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__183_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__183_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__183_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__183_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__183_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__183_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__183_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__183_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__183_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__183_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__183_ccff_tail));

	tile_1__2_ tile_17__16_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_18__2__8_cbx_18__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__6__17_cby_1__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_185_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__173_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__185_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[28]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__184_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__184_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__184_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__184_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__184_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__184_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__184_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__184_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__184_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__184_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__184_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__184_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__184_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__184_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__184_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__184_ccff_tail));

	tile_1__2_ tile_17__17_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__184_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__184_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__184_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__184_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__184_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_18__2__9_cbx_18__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__184_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_186_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__174_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__186_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_18__2__9_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__185_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__185_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__185_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__185_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__185_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__185_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__185_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__185_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__185_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__185_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__185_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__185_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__185_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__185_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__185_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__185_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__185_ccff_tail));

	tile_1__2_ tile_17__18_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__185_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__185_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__185_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__185_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__185_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_18__2__10_cbx_18__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__185_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__19__16_cbx_1__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_17__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__1__chanx_left_in(tile_1__2__175_sb_1__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__19__16_sb_1__18__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__175_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__186_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__186_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__186_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__186_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__186_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__186_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__186_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__186_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__186_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__186_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__186_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__186_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__186_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__186_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__186_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__186_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__186_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__186_ccff_tail));

	tile_1__5_ tile_1__5_ (
		.prog_clk(prog_clk),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__chany_bottom_in(tile_1__2__2_cby_1__2__chany_top_out[0:64]),
		.sb_2__4__chanx_right_in(tile_1__5__2_cbx_1__4__chanx_left_out[0:64]),
		.sb_2__4__chany_bottom_in(tile_1__2__13_cby_1__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__4__chanx_left_in(tile_0__5__0_sb_0__4__chanx_right_out[0:64]),
		.cby_2__5__chany_top_in(tile_2__6__0_sb_2__5__chany_bottom_out[0:64]),
		.ccff_head(tile_1__5__2_ccff_tail),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__0_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__0_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__4__chany_bottom_out(tile_1__5__0_sb_1__4__chany_bottom_out[0:64]),
		.sb_2__4__chanx_right_out(tile_1__5__0_sb_2__4__chanx_right_out[0:64]),
		.sb_2__4__chany_bottom_out(tile_1__5__0_sb_2__4__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_1__4__chanx_left_out(tile_1__5__0_cbx_1__4__chanx_left_out[0:64]),
		.cby_2__5__chany_top_out(tile_1__5__0_cby_2__5__chany_top_out[0:64]),
		.ccff_tail(tile_1__5__0_ccff_tail));

	tile_1__5_ tile_1__14_ (
		.prog_clk(prog_clk),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__18_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__18_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__18_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__18_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__18_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__chany_bottom_in(tile_1__2__7_cby_1__2__chany_top_out[0:64]),
		.sb_2__4__chanx_right_in(tile_1__5__3_cbx_1__4__chanx_left_out[0:64]),
		.sb_2__4__chany_bottom_in(tile_1__2__18_cby_1__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__4__chanx_left_in(tile_0__5__1_sb_0__4__chanx_right_out[0:64]),
		.cby_2__5__chany_top_in(tile_2__6__1_sb_2__5__chany_bottom_out[0:64]),
		.ccff_head(tile_0__5__1_ccff_tail),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__1_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__1_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__4__chany_bottom_out(tile_1__5__1_sb_1__4__chany_bottom_out[0:64]),
		.sb_2__4__chanx_right_out(tile_1__5__1_sb_2__4__chanx_right_out[0:64]),
		.sb_2__4__chany_bottom_out(tile_1__5__1_sb_2__4__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_1__4__chanx_left_out(tile_1__5__1_cbx_1__4__chanx_left_out[0:64]),
		.cby_2__5__chany_top_out(tile_1__5__1_cby_2__5__chany_top_out[0:64]),
		.ccff_tail(tile_1__5__1_ccff_tail));

	tile_1__5_ tile_3__5_ (
		.prog_clk(prog_clk),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__24_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__24_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__24_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__24_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__24_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__35_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__35_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__35_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__35_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__35_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__chany_bottom_in(tile_1__2__24_cby_1__2__chany_top_out[0:64]),
		.sb_2__4__chanx_right_in(tile_1__5__4_cbx_1__4__chanx_left_out[0:64]),
		.sb_2__4__chany_bottom_in(tile_1__2__35_cby_1__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__4__chanx_left_in(tile_1__5__0_sb_2__4__chanx_right_out[0:64]),
		.cby_2__5__chany_top_in(tile_2__6__2_sb_2__5__chany_bottom_out[0:64]),
		.ccff_head(tile_1__5__4_ccff_tail),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__2_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__2_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__4__chany_bottom_out(tile_1__5__2_sb_1__4__chany_bottom_out[0:64]),
		.sb_2__4__chanx_right_out(tile_1__5__2_sb_2__4__chanx_right_out[0:64]),
		.sb_2__4__chany_bottom_out(tile_1__5__2_sb_2__4__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_1__4__chanx_left_out(tile_1__5__2_cbx_1__4__chanx_left_out[0:64]),
		.cby_2__5__chany_top_out(tile_1__5__2_cby_2__5__chany_top_out[0:64]),
		.ccff_tail(tile_1__5__2_ccff_tail));

	tile_1__5_ tile_3__14_ (
		.prog_clk(prog_clk),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__29_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__29_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__29_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__29_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__29_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__40_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__40_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__40_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__40_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__40_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__chany_bottom_in(tile_1__2__29_cby_1__2__chany_top_out[0:64]),
		.sb_2__4__chanx_right_in(tile_1__5__5_cbx_1__4__chanx_left_out[0:64]),
		.sb_2__4__chany_bottom_in(tile_1__2__40_cby_1__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__4__chanx_left_in(tile_1__5__1_sb_2__4__chanx_right_out[0:64]),
		.cby_2__5__chany_top_in(tile_2__6__3_sb_2__5__chany_bottom_out[0:64]),
		.ccff_head(tile_1__5__1_ccff_tail),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__3_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__3_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__4__chany_bottom_out(tile_1__5__3_sb_1__4__chany_bottom_out[0:64]),
		.sb_2__4__chanx_right_out(tile_1__5__3_sb_2__4__chanx_right_out[0:64]),
		.sb_2__4__chany_bottom_out(tile_1__5__3_sb_2__4__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_1__4__chanx_left_out(tile_1__5__3_cbx_1__4__chanx_left_out[0:64]),
		.cby_2__5__chany_top_out(tile_1__5__3_cby_2__5__chany_top_out[0:64]),
		.ccff_tail(tile_1__5__3_ccff_tail));

	tile_1__5_ tile_5__5_ (
		.prog_clk(prog_clk),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__46_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__46_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__46_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__46_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__46_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__57_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__57_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__57_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__57_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__57_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__chany_bottom_in(tile_1__2__46_cby_1__2__chany_top_out[0:64]),
		.sb_2__4__chanx_right_in(tile_1__5__6_cbx_1__4__chanx_left_out[0:64]),
		.sb_2__4__chany_bottom_in(tile_1__2__57_cby_1__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__4__chanx_left_in(tile_1__5__2_sb_2__4__chanx_right_out[0:64]),
		.cby_2__5__chany_top_in(tile_2__6__4_sb_2__5__chany_bottom_out[0:64]),
		.ccff_head(tile_1__5__6_ccff_tail),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__4_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__4_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__4__chany_bottom_out(tile_1__5__4_sb_1__4__chany_bottom_out[0:64]),
		.sb_2__4__chanx_right_out(tile_1__5__4_sb_2__4__chanx_right_out[0:64]),
		.sb_2__4__chany_bottom_out(tile_1__5__4_sb_2__4__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_1__4__chanx_left_out(tile_1__5__4_cbx_1__4__chanx_left_out[0:64]),
		.cby_2__5__chany_top_out(tile_1__5__4_cby_2__5__chany_top_out[0:64]),
		.ccff_tail(tile_1__5__4_ccff_tail));

	tile_1__5_ tile_5__14_ (
		.prog_clk(prog_clk),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__51_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__51_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__51_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__51_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__51_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__62_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__62_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__62_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__62_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__62_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__chany_bottom_in(tile_1__2__51_cby_1__2__chany_top_out[0:64]),
		.sb_2__4__chanx_right_in(tile_1__5__7_cbx_1__4__chanx_left_out[0:64]),
		.sb_2__4__chany_bottom_in(tile_1__2__62_cby_1__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__4__chanx_left_in(tile_1__5__3_sb_2__4__chanx_right_out[0:64]),
		.cby_2__5__chany_top_in(tile_2__6__5_sb_2__5__chany_bottom_out[0:64]),
		.ccff_head(tile_1__5__3_ccff_tail),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__5_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__5_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__4__chany_bottom_out(tile_1__5__5_sb_1__4__chany_bottom_out[0:64]),
		.sb_2__4__chanx_right_out(tile_1__5__5_sb_2__4__chanx_right_out[0:64]),
		.sb_2__4__chany_bottom_out(tile_1__5__5_sb_2__4__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_1__4__chanx_left_out(tile_1__5__5_cbx_1__4__chanx_left_out[0:64]),
		.cby_2__5__chany_top_out(tile_1__5__5_cby_2__5__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[23]));

	tile_1__5_ tile_7__5_ (
		.prog_clk(prog_clk),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__68_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__68_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__68_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__68_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__68_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__79_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__79_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__79_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__79_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__79_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__chany_bottom_in(tile_1__2__68_cby_1__2__chany_top_out[0:64]),
		.sb_2__4__chanx_right_in(tile_1__5__8_cbx_1__4__chanx_left_out[0:64]),
		.sb_2__4__chany_bottom_in(tile_1__2__79_cby_1__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__4__chanx_left_in(tile_1__5__4_sb_2__4__chanx_right_out[0:64]),
		.cby_2__5__chany_top_in(tile_2__6__6_sb_2__5__chany_bottom_out[0:64]),
		.ccff_head(tile_1__5__8_ccff_tail),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__6_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__6_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__4__chany_bottom_out(tile_1__5__6_sb_1__4__chany_bottom_out[0:64]),
		.sb_2__4__chanx_right_out(tile_1__5__6_sb_2__4__chanx_right_out[0:64]),
		.sb_2__4__chany_bottom_out(tile_1__5__6_sb_2__4__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_1__4__chanx_left_out(tile_1__5__6_cbx_1__4__chanx_left_out[0:64]),
		.cby_2__5__chany_top_out(tile_1__5__6_cby_2__5__chany_top_out[0:64]),
		.ccff_tail(tile_1__5__6_ccff_tail));

	tile_1__5_ tile_7__14_ (
		.prog_clk(prog_clk),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__73_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__73_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__73_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__73_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__73_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__84_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__84_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__84_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__84_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__84_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__chany_bottom_in(tile_1__2__73_cby_1__2__chany_top_out[0:64]),
		.sb_2__4__chanx_right_in(tile_1__5__9_cbx_1__4__chanx_left_out[0:64]),
		.sb_2__4__chany_bottom_in(tile_1__2__84_cby_1__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__4__chanx_left_in(tile_1__5__5_sb_2__4__chanx_right_out[0:64]),
		.cby_2__5__chany_top_in(tile_2__6__7_sb_2__5__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[24]),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__7_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__7_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__4__chany_bottom_out(tile_1__5__7_sb_1__4__chany_bottom_out[0:64]),
		.sb_2__4__chanx_right_out(tile_1__5__7_sb_2__4__chanx_right_out[0:64]),
		.sb_2__4__chany_bottom_out(tile_1__5__7_sb_2__4__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_1__4__chanx_left_out(tile_1__5__7_cbx_1__4__chanx_left_out[0:64]),
		.cby_2__5__chany_top_out(tile_1__5__7_cby_2__5__chany_top_out[0:64]),
		.ccff_tail(tile_1__5__7_ccff_tail));

	tile_1__5_ tile_9__5_ (
		.prog_clk(prog_clk),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__90_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__90_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__90_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__90_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__90_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__101_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__101_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__101_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__101_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__101_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__chany_bottom_in(tile_1__2__90_cby_1__2__chany_top_out[0:64]),
		.sb_2__4__chanx_right_in(tile_1__5__10_cbx_1__4__chanx_left_out[0:64]),
		.sb_2__4__chany_bottom_in(tile_1__2__101_cby_1__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__4__chanx_left_in(tile_1__5__6_sb_2__4__chanx_right_out[0:64]),
		.cby_2__5__chany_top_in(tile_2__6__8_sb_2__5__chany_bottom_out[0:64]),
		.ccff_head(tile_1__5__10_ccff_tail),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__8_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__8_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__4__chany_bottom_out(tile_1__5__8_sb_1__4__chany_bottom_out[0:64]),
		.sb_2__4__chanx_right_out(tile_1__5__8_sb_2__4__chanx_right_out[0:64]),
		.sb_2__4__chany_bottom_out(tile_1__5__8_sb_2__4__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_1__4__chanx_left_out(tile_1__5__8_cbx_1__4__chanx_left_out[0:64]),
		.cby_2__5__chany_top_out(tile_1__5__8_cby_2__5__chany_top_out[0:64]),
		.ccff_tail(tile_1__5__8_ccff_tail));

	tile_1__5_ tile_9__14_ (
		.prog_clk(prog_clk),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__95_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__95_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__95_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__95_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__95_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__106_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__106_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__106_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__106_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__106_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__chany_bottom_in(tile_1__2__95_cby_1__2__chany_top_out[0:64]),
		.sb_2__4__chanx_right_in(tile_1__5__11_cbx_1__4__chanx_left_out[0:64]),
		.sb_2__4__chany_bottom_in(tile_1__2__106_cby_1__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__4__chanx_left_in(tile_1__5__7_sb_2__4__chanx_right_out[0:64]),
		.cby_2__5__chany_top_in(tile_2__6__9_sb_2__5__chany_bottom_out[0:64]),
		.ccff_head(tile_1__5__7_ccff_tail),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__9_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__9_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__4__chany_bottom_out(tile_1__5__9_sb_1__4__chany_bottom_out[0:64]),
		.sb_2__4__chanx_right_out(tile_1__5__9_sb_2__4__chanx_right_out[0:64]),
		.sb_2__4__chany_bottom_out(tile_1__5__9_sb_2__4__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_1__4__chanx_left_out(tile_1__5__9_cbx_1__4__chanx_left_out[0:64]),
		.cby_2__5__chany_top_out(tile_1__5__9_cby_2__5__chany_top_out[0:64]),
		.ccff_tail(tile_1__5__9_ccff_tail));

	tile_1__5_ tile_11__5_ (
		.prog_clk(prog_clk),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__112_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__112_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__112_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__112_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__112_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__123_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__123_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__123_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__123_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__123_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__chany_bottom_in(tile_1__2__112_cby_1__2__chany_top_out[0:64]),
		.sb_2__4__chanx_right_in(tile_1__5__12_cbx_1__4__chanx_left_out[0:64]),
		.sb_2__4__chany_bottom_in(tile_1__2__123_cby_1__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__4__chanx_left_in(tile_1__5__8_sb_2__4__chanx_right_out[0:64]),
		.cby_2__5__chany_top_in(tile_2__6__10_sb_2__5__chany_bottom_out[0:64]),
		.ccff_head(tile_1__5__12_ccff_tail),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__10_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__10_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__4__chany_bottom_out(tile_1__5__10_sb_1__4__chany_bottom_out[0:64]),
		.sb_2__4__chanx_right_out(tile_1__5__10_sb_2__4__chanx_right_out[0:64]),
		.sb_2__4__chany_bottom_out(tile_1__5__10_sb_2__4__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_1__4__chanx_left_out(tile_1__5__10_cbx_1__4__chanx_left_out[0:64]),
		.cby_2__5__chany_top_out(tile_1__5__10_cby_2__5__chany_top_out[0:64]),
		.ccff_tail(tile_1__5__10_ccff_tail));

	tile_1__5_ tile_11__14_ (
		.prog_clk(prog_clk),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__117_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__117_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__117_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__117_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__117_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__128_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__128_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__128_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__128_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__128_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__chany_bottom_in(tile_1__2__117_cby_1__2__chany_top_out[0:64]),
		.sb_2__4__chanx_right_in(tile_1__5__13_cbx_1__4__chanx_left_out[0:64]),
		.sb_2__4__chany_bottom_in(tile_1__2__128_cby_1__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__4__chanx_left_in(tile_1__5__9_sb_2__4__chanx_right_out[0:64]),
		.cby_2__5__chany_top_in(tile_2__6__11_sb_2__5__chany_bottom_out[0:64]),
		.ccff_head(tile_1__5__9_ccff_tail),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__11_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__11_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__4__chany_bottom_out(tile_1__5__11_sb_1__4__chany_bottom_out[0:64]),
		.sb_2__4__chanx_right_out(tile_1__5__11_sb_2__4__chanx_right_out[0:64]),
		.sb_2__4__chany_bottom_out(tile_1__5__11_sb_2__4__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_1__4__chanx_left_out(tile_1__5__11_cbx_1__4__chanx_left_out[0:64]),
		.cby_2__5__chany_top_out(tile_1__5__11_cby_2__5__chany_top_out[0:64]),
		.ccff_tail(tile_1__5__11_ccff_tail));

	tile_1__5_ tile_13__5_ (
		.prog_clk(prog_clk),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__134_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__134_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__134_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__134_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__134_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__145_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__145_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__145_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__145_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__145_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__chany_bottom_in(tile_1__2__134_cby_1__2__chany_top_out[0:64]),
		.sb_2__4__chanx_right_in(tile_1__5__14_cbx_1__4__chanx_left_out[0:64]),
		.sb_2__4__chany_bottom_in(tile_1__2__145_cby_1__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__4__chanx_left_in(tile_1__5__10_sb_2__4__chanx_right_out[0:64]),
		.cby_2__5__chany_top_in(tile_2__6__12_sb_2__5__chany_bottom_out[0:64]),
		.ccff_head(tile_1__5__14_ccff_tail),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__12_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__12_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__4__chany_bottom_out(tile_1__5__12_sb_1__4__chany_bottom_out[0:64]),
		.sb_2__4__chanx_right_out(tile_1__5__12_sb_2__4__chanx_right_out[0:64]),
		.sb_2__4__chany_bottom_out(tile_1__5__12_sb_2__4__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_1__4__chanx_left_out(tile_1__5__12_cbx_1__4__chanx_left_out[0:64]),
		.cby_2__5__chany_top_out(tile_1__5__12_cby_2__5__chany_top_out[0:64]),
		.ccff_tail(tile_1__5__12_ccff_tail));

	tile_1__5_ tile_13__14_ (
		.prog_clk(prog_clk),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__139_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__139_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__139_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__139_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__139_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__150_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__150_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__150_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__150_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__150_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__chany_bottom_in(tile_1__2__139_cby_1__2__chany_top_out[0:64]),
		.sb_2__4__chanx_right_in(tile_1__5__15_cbx_1__4__chanx_left_out[0:64]),
		.sb_2__4__chany_bottom_in(tile_1__2__150_cby_1__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__4__chanx_left_in(tile_1__5__11_sb_2__4__chanx_right_out[0:64]),
		.cby_2__5__chany_top_in(tile_2__6__13_sb_2__5__chany_bottom_out[0:64]),
		.ccff_head(tile_1__5__11_ccff_tail),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__13_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__13_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__4__chany_bottom_out(tile_1__5__13_sb_1__4__chany_bottom_out[0:64]),
		.sb_2__4__chanx_right_out(tile_1__5__13_sb_2__4__chanx_right_out[0:64]),
		.sb_2__4__chany_bottom_out(tile_1__5__13_sb_2__4__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_1__4__chanx_left_out(tile_1__5__13_cbx_1__4__chanx_left_out[0:64]),
		.cby_2__5__chany_top_out(tile_1__5__13_cby_2__5__chany_top_out[0:64]),
		.ccff_tail(tile_1__5__13_ccff_tail));

	tile_1__5_ tile_15__5_ (
		.prog_clk(prog_clk),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__156_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__156_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__156_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__156_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__156_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__167_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__167_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__167_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__167_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__167_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__chany_bottom_in(tile_1__2__156_cby_1__2__chany_top_out[0:64]),
		.sb_2__4__chanx_right_in(tile_17__5__0_cbx_17__4__chanx_left_out[0:64]),
		.sb_2__4__chany_bottom_in(tile_1__2__167_cby_1__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__4__chanx_left_in(tile_1__5__12_sb_2__4__chanx_right_out[0:64]),
		.cby_2__5__chany_top_in(tile_2__6__14_sb_2__5__chany_bottom_out[0:64]),
		.ccff_head(tile_17__5__0_ccff_tail),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__14_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__14_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__4__chany_bottom_out(tile_1__5__14_sb_1__4__chany_bottom_out[0:64]),
		.sb_2__4__chanx_right_out(tile_1__5__14_sb_2__4__chanx_right_out[0:64]),
		.sb_2__4__chany_bottom_out(tile_1__5__14_sb_2__4__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_1__4__chanx_left_out(tile_1__5__14_cbx_1__4__chanx_left_out[0:64]),
		.cby_2__5__chany_top_out(tile_1__5__14_cby_2__5__chany_top_out[0:64]),
		.ccff_tail(tile_1__5__14_ccff_tail));

	tile_1__5_ tile_15__14_ (
		.prog_clk(prog_clk),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__161_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__161_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__161_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__161_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__161_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__172_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__172_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__172_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__172_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__172_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__4__chany_bottom_in(tile_1__2__161_cby_1__2__chany_top_out[0:64]),
		.sb_2__4__chanx_right_in(tile_17__5__1_cbx_17__4__chanx_left_out[0:64]),
		.sb_2__4__chany_bottom_in(tile_1__2__172_cby_1__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__4__chanx_left_in(tile_1__5__13_sb_2__4__chanx_right_out[0:64]),
		.cby_2__5__chany_top_in(tile_2__6__15_sb_2__5__chany_bottom_out[0:64]),
		.ccff_head(tile_1__5__13_ccff_tail),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__15_cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__5__15_cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__4__chany_bottom_out(tile_1__5__15_sb_1__4__chany_bottom_out[0:64]),
		.sb_2__4__chanx_right_out(tile_1__5__15_sb_2__4__chanx_right_out[0:64]),
		.sb_2__4__chany_bottom_out(tile_1__5__15_sb_2__4__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_1__4__chanx_left_out(tile_1__5__15_cbx_1__4__chanx_left_out[0:64]),
		.cby_2__5__chany_top_out(tile_1__5__15_cby_2__5__chany_top_out[0:64]),
		.ccff_tail(tile_1__5__15_ccff_tail));

	tile_1__6_ tile_1__6_ (
		.prog_clk(prog_clk),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_1__5__chanx_right_in(tile_2__6__0_cbx_2__5__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_3_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__5__chanx_left_in(tile_0__6__0_sb_0__5__chanx_right_out[0:64]),
		.cby_1__6__chany_top_in(tile_1__2__3_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[10]),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__0_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.sb_1__5__chanx_right_out(tile_1__6__0_sb_1__5__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__5__chanx_left_out(tile_1__6__0_cbx_1__5__chanx_left_out[0:64]),
		.cby_1__6__chany_top_out(tile_1__6__0_cby_1__6__chany_top_out[0:64]),
		.ccff_tail(tile_1__6__0_ccff_tail));

	tile_1__6_ tile_1__15_ (
		.prog_clk(prog_clk),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_1__5__chanx_right_in(tile_2__6__1_cbx_2__5__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__8_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_8_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__5__chanx_left_in(tile_0__6__1_sb_0__5__chanx_right_out[0:64]),
		.cby_1__6__chany_top_in(tile_1__2__8_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__6__1_ccff_tail),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__1_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.sb_1__5__chanx_right_out(tile_1__6__1_sb_1__5__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__5__chanx_left_out(tile_1__6__1_cbx_1__5__chanx_left_out[0:64]),
		.cby_1__6__chany_top_out(tile_1__6__1_cby_1__6__chany_top_out[0:64]),
		.ccff_tail(tile_1__6__1_ccff_tail));

	tile_1__6_ tile_3__6_ (
		.prog_clk(prog_clk),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_1__5__chanx_right_in(tile_2__6__2_cbx_2__5__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__25_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_25_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__5__chanx_left_in(tile_2__6__0_sb_2__5__chanx_right_out[0:64]),
		.cby_1__6__chany_top_in(tile_1__2__25_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__6__0_ccff_tail),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__2_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.sb_1__5__chanx_right_out(tile_1__6__2_sb_1__5__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_3__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__5__chanx_left_out(tile_1__6__2_cbx_1__5__chanx_left_out[0:64]),
		.cby_1__6__chany_top_out(tile_1__6__2_cby_1__6__chany_top_out[0:64]),
		.ccff_tail(tile_1__6__2_ccff_tail));

	tile_1__6_ tile_3__15_ (
		.prog_clk(prog_clk),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_1__5__chanx_right_in(tile_2__6__3_cbx_2__5__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__30_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_30_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__5__chanx_left_in(tile_2__6__1_sb_2__5__chanx_right_out[0:64]),
		.cby_1__6__chany_top_in(tile_1__2__30_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__6__3_ccff_tail),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__3_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.sb_1__5__chanx_right_out(tile_1__6__3_sb_1__5__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_3__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__5__chanx_left_out(tile_1__6__3_cbx_1__5__chanx_left_out[0:64]),
		.cby_1__6__chany_top_out(tile_1__6__3_cby_1__6__chany_top_out[0:64]),
		.ccff_tail(tile_1__6__3_ccff_tail));

	tile_1__6_ tile_5__6_ (
		.prog_clk(prog_clk),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_1__5__chanx_right_in(tile_2__6__4_cbx_2__5__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__47_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_47_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__5__chanx_left_in(tile_2__6__2_sb_2__5__chanx_right_out[0:64]),
		.cby_1__6__chany_top_in(tile_1__2__47_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__6__2_ccff_tail),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__4_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.sb_1__5__chanx_right_out(tile_1__6__4_sb_1__5__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_5__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__5__chanx_left_out(tile_1__6__4_cbx_1__5__chanx_left_out[0:64]),
		.cby_1__6__chany_top_out(tile_1__6__4_cby_1__6__chany_top_out[0:64]),
		.ccff_tail(tile_1__6__4_ccff_tail));

	tile_1__6_ tile_5__15_ (
		.prog_clk(prog_clk),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_1__5__chanx_right_in(tile_2__6__5_cbx_2__5__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__52_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_52_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__5__chanx_left_in(tile_2__6__3_sb_2__5__chanx_right_out[0:64]),
		.cby_1__6__chany_top_in(tile_1__2__52_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__6__5_ccff_tail),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__5_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.sb_1__5__chanx_right_out(tile_1__6__5_sb_1__5__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_5__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__5__chanx_left_out(tile_1__6__5_cbx_1__5__chanx_left_out[0:64]),
		.cby_1__6__chany_top_out(tile_1__6__5_cby_1__6__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[25]));

	tile_1__6_ tile_7__6_ (
		.prog_clk(prog_clk),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_1__5__chanx_right_in(tile_2__6__6_cbx_2__5__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__69_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_69_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__5__chanx_left_in(tile_2__6__4_sb_2__5__chanx_right_out[0:64]),
		.cby_1__6__chany_top_in(tile_1__2__69_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__6__4_ccff_tail),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__6_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.sb_1__5__chanx_right_out(tile_1__6__6_sb_1__5__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_7__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__5__chanx_left_out(tile_1__6__6_cbx_1__5__chanx_left_out[0:64]),
		.cby_1__6__chany_top_out(tile_1__6__6_cby_1__6__chany_top_out[0:64]),
		.ccff_tail(tile_1__6__6_ccff_tail));

	tile_1__6_ tile_7__15_ (
		.prog_clk(prog_clk),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_1__5__chanx_right_in(tile_2__6__7_cbx_2__5__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__74_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_74_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__5__chanx_left_in(tile_2__6__5_sb_2__5__chanx_right_out[0:64]),
		.cby_1__6__chany_top_in(tile_1__2__74_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__6__7_ccff_tail),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__7_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.sb_1__5__chanx_right_out(tile_1__6__7_sb_1__5__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_7__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__5__chanx_left_out(tile_1__6__7_cbx_1__5__chanx_left_out[0:64]),
		.cby_1__6__chany_top_out(tile_1__6__7_cby_1__6__chany_top_out[0:64]),
		.ccff_tail(tile_1__6__7_ccff_tail));

	tile_1__6_ tile_9__6_ (
		.prog_clk(prog_clk),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_1__5__chanx_right_in(tile_2__6__8_cbx_2__5__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__91_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_91_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__5__chanx_left_in(tile_2__6__6_sb_2__5__chanx_right_out[0:64]),
		.cby_1__6__chany_top_in(tile_1__2__91_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__6__6_ccff_tail),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__8_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.sb_1__5__chanx_right_out(tile_1__6__8_sb_1__5__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_9__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__5__chanx_left_out(tile_1__6__8_cbx_1__5__chanx_left_out[0:64]),
		.cby_1__6__chany_top_out(tile_1__6__8_cby_1__6__chany_top_out[0:64]),
		.ccff_tail(tile_1__6__8_ccff_tail));

	tile_1__6_ tile_9__15_ (
		.prog_clk(prog_clk),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_1__5__chanx_right_in(tile_2__6__9_cbx_2__5__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__96_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_96_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__5__chanx_left_in(tile_2__6__7_sb_2__5__chanx_right_out[0:64]),
		.cby_1__6__chany_top_in(tile_1__2__96_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__6__9_ccff_tail),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__9_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.sb_1__5__chanx_right_out(tile_1__6__9_sb_1__5__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_9__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__5__chanx_left_out(tile_1__6__9_cbx_1__5__chanx_left_out[0:64]),
		.cby_1__6__chany_top_out(tile_1__6__9_cby_1__6__chany_top_out[0:64]),
		.ccff_tail(tile_1__6__9_ccff_tail));

	tile_1__6_ tile_11__6_ (
		.prog_clk(prog_clk),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_1__5__chanx_right_in(tile_2__6__10_cbx_2__5__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__113_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_113_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__5__chanx_left_in(tile_2__6__8_sb_2__5__chanx_right_out[0:64]),
		.cby_1__6__chany_top_in(tile_1__2__113_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__6__8_ccff_tail),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__10_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.sb_1__5__chanx_right_out(tile_1__6__10_sb_1__5__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_11__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__5__chanx_left_out(tile_1__6__10_cbx_1__5__chanx_left_out[0:64]),
		.cby_1__6__chany_top_out(tile_1__6__10_cby_1__6__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[10]));

	tile_1__6_ tile_11__15_ (
		.prog_clk(prog_clk),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_1__5__chanx_right_in(tile_2__6__11_cbx_2__5__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__118_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_118_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__5__chanx_left_in(tile_2__6__9_sb_2__5__chanx_right_out[0:64]),
		.cby_1__6__chany_top_in(tile_1__2__118_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__6__11_ccff_tail),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__11_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.sb_1__5__chanx_right_out(tile_1__6__11_sb_1__5__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_11__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__5__chanx_left_out(tile_1__6__11_cbx_1__5__chanx_left_out[0:64]),
		.cby_1__6__chany_top_out(tile_1__6__11_cby_1__6__chany_top_out[0:64]),
		.ccff_tail(tile_1__6__11_ccff_tail));

	tile_1__6_ tile_13__6_ (
		.prog_clk(prog_clk),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_1__5__chanx_right_in(tile_2__6__12_cbx_2__5__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__135_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_135_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__5__chanx_left_in(tile_2__6__10_sb_2__5__chanx_right_out[0:64]),
		.cby_1__6__chany_top_in(tile_1__2__135_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__6__10_ccff_tail),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__12_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.sb_1__5__chanx_right_out(tile_1__6__12_sb_1__5__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_13__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__5__chanx_left_out(tile_1__6__12_cbx_1__5__chanx_left_out[0:64]),
		.cby_1__6__chany_top_out(tile_1__6__12_cby_1__6__chany_top_out[0:64]),
		.ccff_tail(tile_1__6__12_ccff_tail));

	tile_1__6_ tile_13__15_ (
		.prog_clk(prog_clk),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_1__5__chanx_right_in(tile_2__6__13_cbx_2__5__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__140_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_140_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__5__chanx_left_in(tile_2__6__11_sb_2__5__chanx_right_out[0:64]),
		.cby_1__6__chany_top_in(tile_1__2__140_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__6__13_ccff_tail),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__13_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.sb_1__5__chanx_right_out(tile_1__6__13_sb_1__5__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_13__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__5__chanx_left_out(tile_1__6__13_cbx_1__5__chanx_left_out[0:64]),
		.cby_1__6__chany_top_out(tile_1__6__13_cby_1__6__chany_top_out[0:64]),
		.ccff_tail(tile_1__6__13_ccff_tail));

	tile_1__6_ tile_15__6_ (
		.prog_clk(prog_clk),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_1__5__chanx_right_in(tile_2__6__14_cbx_2__5__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__157_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_157_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__5__chanx_left_in(tile_2__6__12_sb_2__5__chanx_right_out[0:64]),
		.cby_1__6__chany_top_in(tile_1__2__157_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__6__12_ccff_tail),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__14_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.sb_1__5__chanx_right_out(tile_1__6__14_sb_1__5__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_15__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__5__chanx_left_out(tile_1__6__14_cbx_1__5__chanx_left_out[0:64]),
		.cby_1__6__chany_top_out(tile_1__6__14_cby_1__6__chany_top_out[0:64]),
		.ccff_tail(tile_1__6__14_ccff_tail));

	tile_1__6_ tile_15__15_ (
		.prog_clk(prog_clk),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_1__5__chanx_right_in(tile_2__6__15_cbx_2__5__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__162_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_162_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__5__chanx_left_in(tile_2__6__13_sb_2__5__chanx_right_out[0:64]),
		.cby_1__6__chany_top_in(tile_1__2__162_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[25]),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__15_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.sb_1__5__chanx_right_out(tile_1__6__15_sb_1__5__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_15__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__5__chanx_left_out(tile_1__6__15_cbx_1__5__chanx_left_out[0:64]),
		.cby_1__6__chany_top_out(tile_1__6__15_cby_1__6__chany_top_out[0:64]),
		.ccff_tail(tile_1__6__15_ccff_tail));

	tile_1__6_ tile_17__6_ (
		.prog_clk(prog_clk),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_1__5__chanx_right_in(tile_18__6__0_cbx_18__5__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__179_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_179_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__5__chanx_left_in(tile_2__6__14_sb_2__5__chanx_right_out[0:64]),
		.cby_1__6__chany_top_in(tile_1__2__179_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__6__14_ccff_tail),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.sb_1__5__chanx_right_out(tile_1__6__16_sb_1__5__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_17__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__5__chanx_left_out(tile_1__6__16_cbx_1__5__chanx_left_out[0:64]),
		.cby_1__6__chany_top_out(tile_1__6__16_cby_1__6__chany_top_out[0:64]),
		.ccff_tail(tile_1__6__16_ccff_tail));

	tile_1__6_ tile_17__15_ (
		.prog_clk(prog_clk),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_1__5__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_1__5__chanx_right_in(tile_18__6__2_cbx_18__5__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__184_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_184_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__5__chanx_left_in(tile_2__6__15_sb_2__5__chanx_right_out[0:64]),
		.cby_1__6__chany_top_in(tile_1__2__184_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_18__6__2_ccff_tail),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.sb_1__5__chanx_right_out(tile_1__6__17_sb_1__5__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__6__17_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__6__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__6__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__6__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__6__17_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_17__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__5__chanx_left_out(tile_1__6__17_cbx_1__5__chanx_left_out[0:64]),
		.cby_1__6__chany_top_out(tile_1__6__17_cby_1__6__chany_top_out[0:64]),
		.ccff_tail(tile_1__6__17_ccff_tail));

	tile_1__10_ tile_1__10_ (
		.prog_clk(prog_clk),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__16_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__16_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__9__chany_bottom_in(tile_1__2__5_cby_1__2__chany_top_out[0:64]),
		.sb_2__9__chanx_right_in(tile_1__10__1_cbx_1__9__chanx_left_out[0:64]),
		.sb_2__9__chany_bottom_in(tile_1__2__16_cby_1__2__chany_top_out[0:64]),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.cbx_1__9__chanx_left_in(tile_0__10__0_sb_0__9__chanx_right_out[0:64]),
		.cby_2__10__chany_top_in(tile_2__11__0_sb_2__10__chany_bottom_out[0:64]),
		.ccff_head(tile_0__10__0_ccff_tail),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__0_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__0_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__9__chany_bottom_out(tile_1__10__0_sb_1__9__chany_bottom_out[0:64]),
		.sb_2__9__chanx_right_out(tile_1__10__0_sb_2__9__chanx_right_out[0:64]),
		.sb_2__9__chany_bottom_out(tile_1__10__0_sb_2__9__chany_bottom_out[0:64]),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_1__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.cbx_1__9__chanx_left_out(tile_1__10__0_cbx_1__9__chanx_left_out[0:64]),
		.cby_2__10__chany_top_out(tile_1__10__0_cby_2__10__chany_top_out[0:64]),
		.ccff_tail(tile_1__10__0_ccff_tail));

	tile_1__10_ tile_3__10_ (
		.prog_clk(prog_clk),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__27_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__27_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__27_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__27_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__27_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__38_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__38_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__38_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__38_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__38_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__9__chany_bottom_in(tile_1__2__27_cby_1__2__chany_top_out[0:64]),
		.sb_2__9__chanx_right_in(tile_1__10__2_cbx_1__9__chanx_left_out[0:64]),
		.sb_2__9__chany_bottom_in(tile_1__2__38_cby_1__2__chany_top_out[0:64]),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.cbx_1__9__chanx_left_in(tile_1__10__0_sb_2__9__chanx_right_out[0:64]),
		.cby_2__10__chany_top_in(tile_2__11__1_sb_2__10__chany_bottom_out[0:64]),
		.ccff_head(tile_1__10__0_ccff_tail),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__1_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__1_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__9__chany_bottom_out(tile_1__10__1_sb_1__9__chany_bottom_out[0:64]),
		.sb_2__9__chanx_right_out(tile_1__10__1_sb_2__9__chanx_right_out[0:64]),
		.sb_2__9__chany_bottom_out(tile_1__10__1_sb_2__9__chany_bottom_out[0:64]),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_1__10__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.cbx_1__9__chanx_left_out(tile_1__10__1_cbx_1__9__chanx_left_out[0:64]),
		.cby_2__10__chany_top_out(tile_1__10__1_cby_2__10__chany_top_out[0:64]),
		.ccff_tail(tile_1__10__1_ccff_tail));

	tile_1__10_ tile_5__10_ (
		.prog_clk(prog_clk),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__49_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__49_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__49_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__49_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__49_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__60_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__60_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__60_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__60_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__60_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__9__chany_bottom_in(tile_1__2__49_cby_1__2__chany_top_out[0:64]),
		.sb_2__9__chanx_right_in(tile_1__10__3_cbx_1__9__chanx_left_out[0:64]),
		.sb_2__9__chany_bottom_in(tile_1__2__60_cby_1__2__chany_top_out[0:64]),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.cbx_1__9__chanx_left_in(tile_1__10__1_sb_2__9__chanx_right_out[0:64]),
		.cby_2__10__chany_top_in(tile_2__11__2_sb_2__10__chany_bottom_out[0:64]),
		.ccff_head(tile_1__10__1_ccff_tail),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__2_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__2_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__9__chany_bottom_out(tile_1__10__2_sb_1__9__chany_bottom_out[0:64]),
		.sb_2__9__chanx_right_out(tile_1__10__2_sb_2__9__chanx_right_out[0:64]),
		.sb_2__9__chany_bottom_out(tile_1__10__2_sb_2__9__chany_bottom_out[0:64]),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_1__10__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.cbx_1__9__chanx_left_out(tile_1__10__2_cbx_1__9__chanx_left_out[0:64]),
		.cby_2__10__chany_top_out(tile_1__10__2_cby_2__10__chany_top_out[0:64]),
		.ccff_tail(tile_1__10__2_ccff_tail));

	tile_1__10_ tile_7__10_ (
		.prog_clk(prog_clk),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__71_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__71_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__71_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__71_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__71_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__82_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__82_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__82_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__82_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__82_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__9__chany_bottom_in(tile_1__2__71_cby_1__2__chany_top_out[0:64]),
		.sb_2__9__chanx_right_in(tile_1__10__4_cbx_1__9__chanx_left_out[0:64]),
		.sb_2__9__chany_bottom_in(tile_1__2__82_cby_1__2__chany_top_out[0:64]),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.cbx_1__9__chanx_left_in(tile_1__10__2_sb_2__9__chanx_right_out[0:64]),
		.cby_2__10__chany_top_in(tile_2__11__3_sb_2__10__chany_bottom_out[0:64]),
		.ccff_head(tile_1__10__2_ccff_tail),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__3_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__3_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__9__chany_bottom_out(tile_1__10__3_sb_1__9__chany_bottom_out[0:64]),
		.sb_2__9__chanx_right_out(tile_1__10__3_sb_2__9__chanx_right_out[0:64]),
		.sb_2__9__chany_bottom_out(tile_1__10__3_sb_2__9__chany_bottom_out[0:64]),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_1__10__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.cbx_1__9__chanx_left_out(tile_1__10__3_cbx_1__9__chanx_left_out[0:64]),
		.cby_2__10__chany_top_out(tile_1__10__3_cby_2__10__chany_top_out[0:64]),
		.ccff_tail(tile_1__10__3_ccff_tail));

	tile_1__10_ tile_9__10_ (
		.prog_clk(prog_clk),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__93_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__93_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__93_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__93_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__93_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__104_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__104_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__104_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__104_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__104_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__9__chany_bottom_in(tile_1__2__93_cby_1__2__chany_top_out[0:64]),
		.sb_2__9__chanx_right_in(tile_1__10__5_cbx_1__9__chanx_left_out[0:64]),
		.sb_2__9__chany_bottom_in(tile_1__2__104_cby_1__2__chany_top_out[0:64]),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.cbx_1__9__chanx_left_in(tile_1__10__3_sb_2__9__chanx_right_out[0:64]),
		.cby_2__10__chany_top_in(tile_2__11__4_sb_2__10__chany_bottom_out[0:64]),
		.ccff_head(tile_1__10__3_ccff_tail),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__4_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__4_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__9__chany_bottom_out(tile_1__10__4_sb_1__9__chany_bottom_out[0:64]),
		.sb_2__9__chanx_right_out(tile_1__10__4_sb_2__9__chanx_right_out[0:64]),
		.sb_2__9__chany_bottom_out(tile_1__10__4_sb_2__9__chany_bottom_out[0:64]),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_1__10__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.cbx_1__9__chanx_left_out(tile_1__10__4_cbx_1__9__chanx_left_out[0:64]),
		.cby_2__10__chany_top_out(tile_1__10__4_cby_2__10__chany_top_out[0:64]),
		.ccff_tail(tile_1__10__4_ccff_tail));

	tile_1__10_ tile_11__10_ (
		.prog_clk(prog_clk),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__115_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__115_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__115_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__115_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__115_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__126_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__126_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__126_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__126_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__126_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__9__chany_bottom_in(tile_1__2__115_cby_1__2__chany_top_out[0:64]),
		.sb_2__9__chanx_right_in(tile_1__10__6_cbx_1__9__chanx_left_out[0:64]),
		.sb_2__9__chany_bottom_in(tile_1__2__126_cby_1__2__chany_top_out[0:64]),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.cbx_1__9__chanx_left_in(tile_1__10__4_sb_2__9__chanx_right_out[0:64]),
		.cby_2__10__chany_top_in(tile_2__11__5_sb_2__10__chany_bottom_out[0:64]),
		.ccff_head(tile_1__10__4_ccff_tail),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__5_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__5_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__9__chany_bottom_out(tile_1__10__5_sb_1__9__chany_bottom_out[0:64]),
		.sb_2__9__chanx_right_out(tile_1__10__5_sb_2__9__chanx_right_out[0:64]),
		.sb_2__9__chany_bottom_out(tile_1__10__5_sb_2__9__chany_bottom_out[0:64]),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_1__10__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.cbx_1__9__chanx_left_out(tile_1__10__5_cbx_1__9__chanx_left_out[0:64]),
		.cby_2__10__chany_top_out(tile_1__10__5_cby_2__10__chany_top_out[0:64]),
		.ccff_tail(tile_1__10__5_ccff_tail));

	tile_1__10_ tile_13__10_ (
		.prog_clk(prog_clk),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__137_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__137_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__137_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__137_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__137_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__148_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__148_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__148_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__148_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__148_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__9__chany_bottom_in(tile_1__2__137_cby_1__2__chany_top_out[0:64]),
		.sb_2__9__chanx_right_in(tile_1__10__7_cbx_1__9__chanx_left_out[0:64]),
		.sb_2__9__chany_bottom_in(tile_1__2__148_cby_1__2__chany_top_out[0:64]),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.cbx_1__9__chanx_left_in(tile_1__10__5_sb_2__9__chanx_right_out[0:64]),
		.cby_2__10__chany_top_in(tile_2__11__6_sb_2__10__chany_bottom_out[0:64]),
		.ccff_head(tile_1__10__5_ccff_tail),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__6_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__6_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__9__chany_bottom_out(tile_1__10__6_sb_1__9__chany_bottom_out[0:64]),
		.sb_2__9__chanx_right_out(tile_1__10__6_sb_2__9__chanx_right_out[0:64]),
		.sb_2__9__chany_bottom_out(tile_1__10__6_sb_2__9__chany_bottom_out[0:64]),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_1__10__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.cbx_1__9__chanx_left_out(tile_1__10__6_cbx_1__9__chanx_left_out[0:64]),
		.cby_2__10__chany_top_out(tile_1__10__6_cby_2__10__chany_top_out[0:64]),
		.ccff_tail(tile_1__10__6_ccff_tail));

	tile_1__10_ tile_15__10_ (
		.prog_clk(prog_clk),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__159_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__159_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__159_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__159_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__159_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.sb_2__9__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__170_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__170_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__170_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_2__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__170_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_2__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__170_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__9__chany_bottom_in(tile_1__2__159_cby_1__2__chany_top_out[0:64]),
		.sb_2__9__chanx_right_in(tile_17__10__0_cbx_17__9__chanx_left_out[0:64]),
		.sb_2__9__chany_bottom_in(tile_1__2__170_cby_1__2__chany_top_out[0:64]),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.cbx_1__9__chanx_left_in(tile_1__10__6_sb_2__9__chanx_right_out[0:64]),
		.cby_2__10__chany_top_in(tile_2__11__7_sb_2__10__chany_bottom_out[0:64]),
		.ccff_head(tile_1__10__6_ccff_tail),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__7_cbx_1__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__10__7_cbx_2__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__9__chany_bottom_out(tile_1__10__7_sb_1__9__chany_bottom_out[0:64]),
		.sb_2__9__chanx_right_out(tile_1__10__7_sb_2__9__chanx_right_out[0:64]),
		.sb_2__9__chany_bottom_out(tile_1__10__7_sb_2__9__chany_bottom_out[0:64]),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_1__10__7_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.cbx_1__9__chanx_left_out(tile_1__10__7_cbx_1__9__chanx_left_out[0:64]),
		.cby_2__10__chany_top_out(tile_1__10__7_cby_2__10__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[17]));

	tile_1__11_ tile_1__11_ (
		.prog_clk(prog_clk),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__10__chanx_right_in(tile_2__11__0_cbx_2__10__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_6_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__10__chanx_left_in(tile_0__11__0_sb_0__10__chanx_right_out[0:64]),
		.cby_1__11__chany_top_in(tile_1__2__6_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__11__0_ccff_tail),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_(tile_1__11__0_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.sb_1__10__chanx_right_out(tile_1__11__0_sb_1__10__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__10__chanx_left_out(tile_1__11__0_cbx_1__10__chanx_left_out[0:64]),
		.cby_1__11__chany_top_out(tile_1__11__0_cby_1__11__chany_top_out[0:64]),
		.ccff_tail(tile_1__11__0_ccff_tail));

	tile_1__11_ tile_3__11_ (
		.prog_clk(prog_clk),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__10__chanx_right_in(tile_2__11__1_cbx_2__10__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__28_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_28_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__10__chanx_left_in(tile_2__11__0_sb_2__10__chanx_right_out[0:64]),
		.cby_1__11__chany_top_in(tile_1__2__28_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__11__1_ccff_tail),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_(tile_1__11__1_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.sb_1__10__chanx_right_out(tile_1__11__1_sb_1__10__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_3__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__10__chanx_left_out(tile_1__11__1_cbx_1__10__chanx_left_out[0:64]),
		.cby_1__11__chany_top_out(tile_1__11__1_cby_1__11__chany_top_out[0:64]),
		.ccff_tail(tile_1__11__1_ccff_tail));

	tile_1__11_ tile_5__11_ (
		.prog_clk(prog_clk),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__10__chanx_right_in(tile_2__11__2_cbx_2__10__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__50_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_50_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__10__chanx_left_in(tile_2__11__1_sb_2__10__chanx_right_out[0:64]),
		.cby_1__11__chany_top_in(tile_1__2__50_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__11__2_ccff_tail),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_(tile_1__11__2_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.sb_1__10__chanx_right_out(tile_1__11__2_sb_1__10__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_5__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__10__chanx_left_out(tile_1__11__2_cbx_1__10__chanx_left_out[0:64]),
		.cby_1__11__chany_top_out(tile_1__11__2_cby_1__11__chany_top_out[0:64]),
		.ccff_tail(tile_1__11__2_ccff_tail));

	tile_1__11_ tile_7__11_ (
		.prog_clk(prog_clk),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__10__chanx_right_in(tile_2__11__3_cbx_2__10__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__72_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_72_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__10__chanx_left_in(tile_2__11__2_sb_2__10__chanx_right_out[0:64]),
		.cby_1__11__chany_top_in(tile_1__2__72_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__11__3_ccff_tail),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_(tile_1__11__3_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.sb_1__10__chanx_right_out(tile_1__11__3_sb_1__10__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_7__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__10__chanx_left_out(tile_1__11__3_cbx_1__10__chanx_left_out[0:64]),
		.cby_1__11__chany_top_out(tile_1__11__3_cby_1__11__chany_top_out[0:64]),
		.ccff_tail(tile_1__11__3_ccff_tail));

	tile_1__11_ tile_9__11_ (
		.prog_clk(prog_clk),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__10__chanx_right_in(tile_2__11__4_cbx_2__10__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__94_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_94_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__10__chanx_left_in(tile_2__11__3_sb_2__10__chanx_right_out[0:64]),
		.cby_1__11__chany_top_in(tile_1__2__94_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__11__4_ccff_tail),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_(tile_1__11__4_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.sb_1__10__chanx_right_out(tile_1__11__4_sb_1__10__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_9__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__10__chanx_left_out(tile_1__11__4_cbx_1__10__chanx_left_out[0:64]),
		.cby_1__11__chany_top_out(tile_1__11__4_cby_1__11__chany_top_out[0:64]),
		.ccff_tail(tile_1__11__4_ccff_tail));

	tile_1__11_ tile_11__11_ (
		.prog_clk(prog_clk),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__10__chanx_right_in(tile_2__11__5_cbx_2__10__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__116_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_116_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__10__chanx_left_in(tile_2__11__4_sb_2__10__chanx_right_out[0:64]),
		.cby_1__11__chany_top_in(tile_1__2__116_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__11__5_ccff_tail),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_(tile_1__11__5_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.sb_1__10__chanx_right_out(tile_1__11__5_sb_1__10__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_11__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__10__chanx_left_out(tile_1__11__5_cbx_1__10__chanx_left_out[0:64]),
		.cby_1__11__chany_top_out(tile_1__11__5_cby_1__11__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[18]));

	tile_1__11_ tile_13__11_ (
		.prog_clk(prog_clk),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__10__chanx_right_in(tile_2__11__6_cbx_2__10__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__138_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_138_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__10__chanx_left_in(tile_2__11__5_sb_2__10__chanx_right_out[0:64]),
		.cby_1__11__chany_top_in(tile_1__2__138_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__11__6_ccff_tail),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_(tile_1__11__6_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.sb_1__10__chanx_right_out(tile_1__11__6_sb_1__10__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_13__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__10__chanx_left_out(tile_1__11__6_cbx_1__10__chanx_left_out[0:64]),
		.cby_1__11__chany_top_out(tile_1__11__6_cby_1__11__chany_top_out[0:64]),
		.ccff_tail(tile_1__11__6_ccff_tail));

	tile_1__11_ tile_15__11_ (
		.prog_clk(prog_clk),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__10__chanx_right_in(tile_2__11__7_cbx_2__10__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__160_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_160_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__10__chanx_left_in(tile_2__11__6_sb_2__10__chanx_right_out[0:64]),
		.cby_1__11__chany_top_in(tile_1__2__160_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__11__7_ccff_tail),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_(tile_1__11__7_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.sb_1__10__chanx_right_out(tile_1__11__7_sb_1__10__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_15__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__10__chanx_left_out(tile_1__11__7_cbx_1__10__chanx_left_out[0:64]),
		.cby_1__11__chany_top_out(tile_1__11__7_cby_1__11__chany_top_out[0:64]),
		.ccff_tail(tile_1__11__7_ccff_tail));

	tile_1__11_ tile_17__11_ (
		.prog_clk(prog_clk),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_1__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_1__10__chanx_right_in(tile_18__6__1_cbx_18__5__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__182_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_182_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_1__10__chanx_left_in(tile_2__11__7_sb_2__10__chanx_right_out[0:64]),
		.cby_1__11__chany_top_in(tile_1__2__182_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_18__6__1_ccff_tail),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.sb_1__10__chanx_right_out(tile_1__11__8_sb_1__10__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__11__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__11__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__11__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__11__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__11__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_17__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__11__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__11__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__11__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__11__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__11__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__11__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__10__chanx_left_out(tile_1__11__8_cbx_1__10__chanx_left_out[0:64]),
		.cby_1__11__chany_top_out(tile_1__11__8_cby_1__11__chany_top_out[0:64]),
		.ccff_tail(tile_1__11__8_ccff_tail));

	tile_2__6_ tile_2__6_ (
		.prog_clk(prog_clk),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_2__5__chanx_right_in(tile_1__6__2_cbx_1__5__chanx_left_out[0:64]),
		.sb_2__5__chany_bottom_in(tile_1__5__0_cby_2__5__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__14_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_14_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__5__chanx_left_in(tile_1__6__0_sb_1__5__chanx_right_out[0:64]),
		.cby_2__6__chany_top_in(tile_1__2__14_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__6__0_ccff_tail),
		.sb_2__5__chanx_right_out(tile_2__6__0_sb_2__5__chanx_right_out[0:64]),
		.sb_2__5__chany_bottom_out(tile_2__6__0_sb_2__5__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_2__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__5__chanx_left_out(tile_2__6__0_cbx_2__5__chanx_left_out[0:64]),
		.cby_2__6__chany_top_out(tile_2__6__0_cby_2__6__chany_top_out[0:64]),
		.ccff_tail(tile_2__6__0_ccff_tail));

	tile_2__6_ tile_2__15_ (
		.prog_clk(prog_clk),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_2__5__chanx_right_in(tile_1__6__3_cbx_1__5__chanx_left_out[0:64]),
		.sb_2__5__chany_bottom_in(tile_1__5__1_cby_2__5__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__19_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_19_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__5__chanx_left_in(tile_1__6__1_sb_1__5__chanx_right_out[0:64]),
		.cby_2__6__chany_top_in(tile_1__2__19_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__6__3_ccff_tail),
		.sb_2__5__chanx_right_out(tile_2__6__1_sb_2__5__chanx_right_out[0:64]),
		.sb_2__5__chany_bottom_out(tile_2__6__1_sb_2__5__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_2__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__5__chanx_left_out(tile_2__6__1_cbx_2__5__chanx_left_out[0:64]),
		.cby_2__6__chany_top_out(tile_2__6__1_cby_2__6__chany_top_out[0:64]),
		.ccff_tail(tile_2__6__1_ccff_tail));

	tile_2__6_ tile_4__6_ (
		.prog_clk(prog_clk),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_2__5__chanx_right_in(tile_1__6__4_cbx_1__5__chanx_left_out[0:64]),
		.sb_2__5__chany_bottom_in(tile_1__5__2_cby_2__5__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__36_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_36_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__5__chanx_left_in(tile_1__6__2_sb_1__5__chanx_right_out[0:64]),
		.cby_2__6__chany_top_in(tile_1__2__36_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__6__2_ccff_tail),
		.sb_2__5__chanx_right_out(tile_2__6__2_sb_2__5__chanx_right_out[0:64]),
		.sb_2__5__chany_bottom_out(tile_2__6__2_sb_2__5__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_4__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__5__chanx_left_out(tile_2__6__2_cbx_2__5__chanx_left_out[0:64]),
		.cby_2__6__chany_top_out(tile_2__6__2_cby_2__6__chany_top_out[0:64]),
		.ccff_tail(tile_2__6__2_ccff_tail));

	tile_2__6_ tile_4__15_ (
		.prog_clk(prog_clk),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_2__5__chanx_right_in(tile_1__6__5_cbx_1__5__chanx_left_out[0:64]),
		.sb_2__5__chany_bottom_in(tile_1__5__3_cby_2__5__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__41_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_41_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__5__chanx_left_in(tile_1__6__3_sb_1__5__chanx_right_out[0:64]),
		.cby_2__6__chany_top_in(tile_1__2__41_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[26]),
		.sb_2__5__chanx_right_out(tile_2__6__3_sb_2__5__chanx_right_out[0:64]),
		.sb_2__5__chany_bottom_out(tile_2__6__3_sb_2__5__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_4__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__5__chanx_left_out(tile_2__6__3_cbx_2__5__chanx_left_out[0:64]),
		.cby_2__6__chany_top_out(tile_2__6__3_cby_2__6__chany_top_out[0:64]),
		.ccff_tail(tile_2__6__3_ccff_tail));

	tile_2__6_ tile_6__6_ (
		.prog_clk(prog_clk),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_2__5__chanx_right_in(tile_1__6__6_cbx_1__5__chanx_left_out[0:64]),
		.sb_2__5__chany_bottom_in(tile_1__5__4_cby_2__5__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__58_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_58_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__5__chanx_left_in(tile_1__6__4_sb_1__5__chanx_right_out[0:64]),
		.cby_2__6__chany_top_in(tile_1__2__58_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__6__4_ccff_tail),
		.sb_2__5__chanx_right_out(tile_2__6__4_sb_2__5__chanx_right_out[0:64]),
		.sb_2__5__chany_bottom_out(tile_2__6__4_sb_2__5__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_6__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__5__chanx_left_out(tile_2__6__4_cbx_2__5__chanx_left_out[0:64]),
		.cby_2__6__chany_top_out(tile_2__6__4_cby_2__6__chany_top_out[0:64]),
		.ccff_tail(tile_2__6__4_ccff_tail));

	tile_2__6_ tile_6__15_ (
		.prog_clk(prog_clk),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__7_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_2__5__chanx_right_in(tile_1__6__7_cbx_1__5__chanx_left_out[0:64]),
		.sb_2__5__chany_bottom_in(tile_1__5__5_cby_2__5__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__63_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_63_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__5__chanx_left_in(tile_1__6__5_sb_1__5__chanx_right_out[0:64]),
		.cby_2__6__chany_top_in(tile_1__2__63_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__6__7_ccff_tail),
		.sb_2__5__chanx_right_out(tile_2__6__5_sb_2__5__chanx_right_out[0:64]),
		.sb_2__5__chany_bottom_out(tile_2__6__5_sb_2__5__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_6__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__5__chanx_left_out(tile_2__6__5_cbx_2__5__chanx_left_out[0:64]),
		.cby_2__6__chany_top_out(tile_2__6__5_cby_2__6__chany_top_out[0:64]),
		.ccff_tail(tile_2__6__5_ccff_tail));

	tile_2__6_ tile_8__6_ (
		.prog_clk(prog_clk),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__8_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_2__5__chanx_right_in(tile_1__6__8_cbx_1__5__chanx_left_out[0:64]),
		.sb_2__5__chany_bottom_in(tile_1__5__6_cby_2__5__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__80_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_80_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__5__chanx_left_in(tile_1__6__6_sb_1__5__chanx_right_out[0:64]),
		.cby_2__6__chany_top_in(tile_1__2__80_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__6__6_ccff_tail),
		.sb_2__5__chanx_right_out(tile_2__6__6_sb_2__5__chanx_right_out[0:64]),
		.sb_2__5__chany_bottom_out(tile_2__6__6_sb_2__5__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_8__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__5__chanx_left_out(tile_2__6__6_cbx_2__5__chanx_left_out[0:64]),
		.cby_2__6__chany_top_out(tile_2__6__6_cby_2__6__chany_top_out[0:64]),
		.ccff_tail(tile_2__6__6_ccff_tail));

	tile_2__6_ tile_8__15_ (
		.prog_clk(prog_clk),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__9_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_2__5__chanx_right_in(tile_1__6__9_cbx_1__5__chanx_left_out[0:64]),
		.sb_2__5__chany_bottom_in(tile_1__5__7_cby_2__5__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__85_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_85_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__5__chanx_left_in(tile_1__6__7_sb_1__5__chanx_right_out[0:64]),
		.cby_2__6__chany_top_in(tile_1__2__85_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__6__9_ccff_tail),
		.sb_2__5__chanx_right_out(tile_2__6__7_sb_2__5__chanx_right_out[0:64]),
		.sb_2__5__chany_bottom_out(tile_2__6__7_sb_2__5__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_8__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__5__chanx_left_out(tile_2__6__7_cbx_2__5__chanx_left_out[0:64]),
		.cby_2__6__chany_top_out(tile_2__6__7_cby_2__6__chany_top_out[0:64]),
		.ccff_tail(tile_2__6__7_ccff_tail));

	tile_2__6_ tile_10__6_ (
		.prog_clk(prog_clk),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__10_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_2__5__chanx_right_in(tile_1__6__10_cbx_1__5__chanx_left_out[0:64]),
		.sb_2__5__chany_bottom_in(tile_1__5__8_cby_2__5__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__102_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_102_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__5__chanx_left_in(tile_1__6__8_sb_1__5__chanx_right_out[0:64]),
		.cby_2__6__chany_top_in(tile_1__2__102_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__6__8_ccff_tail),
		.sb_2__5__chanx_right_out(tile_2__6__8_sb_2__5__chanx_right_out[0:64]),
		.sb_2__5__chany_bottom_out(tile_2__6__8_sb_2__5__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_10__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__5__chanx_left_out(tile_2__6__8_cbx_2__5__chanx_left_out[0:64]),
		.cby_2__6__chany_top_out(tile_2__6__8_cby_2__6__chany_top_out[0:64]),
		.ccff_tail(tile_2__6__8_ccff_tail));

	tile_2__6_ tile_10__15_ (
		.prog_clk(prog_clk),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__11_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_2__5__chanx_right_in(tile_1__6__11_cbx_1__5__chanx_left_out[0:64]),
		.sb_2__5__chany_bottom_in(tile_1__5__9_cby_2__5__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__107_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_107_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__5__chanx_left_in(tile_1__6__9_sb_1__5__chanx_right_out[0:64]),
		.cby_2__6__chany_top_in(tile_1__2__107_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__6__11_ccff_tail),
		.sb_2__5__chanx_right_out(tile_2__6__9_sb_2__5__chanx_right_out[0:64]),
		.sb_2__5__chany_bottom_out(tile_2__6__9_sb_2__5__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_10__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__5__chanx_left_out(tile_2__6__9_cbx_2__5__chanx_left_out[0:64]),
		.cby_2__6__chany_top_out(tile_2__6__9_cby_2__6__chany_top_out[0:64]),
		.ccff_tail(tile_2__6__9_ccff_tail));

	tile_2__6_ tile_12__6_ (
		.prog_clk(prog_clk),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__12_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_2__5__chanx_right_in(tile_1__6__12_cbx_1__5__chanx_left_out[0:64]),
		.sb_2__5__chany_bottom_in(tile_1__5__10_cby_2__5__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__124_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_124_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__5__chanx_left_in(tile_1__6__10_sb_1__5__chanx_right_out[0:64]),
		.cby_2__6__chany_top_in(tile_1__2__124_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[11]),
		.sb_2__5__chanx_right_out(tile_2__6__10_sb_2__5__chanx_right_out[0:64]),
		.sb_2__5__chany_bottom_out(tile_2__6__10_sb_2__5__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_12__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__5__chanx_left_out(tile_2__6__10_cbx_2__5__chanx_left_out[0:64]),
		.cby_2__6__chany_top_out(tile_2__6__10_cby_2__6__chany_top_out[0:64]),
		.ccff_tail(tile_2__6__10_ccff_tail));

	tile_2__6_ tile_12__15_ (
		.prog_clk(prog_clk),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__13_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_2__5__chanx_right_in(tile_1__6__13_cbx_1__5__chanx_left_out[0:64]),
		.sb_2__5__chany_bottom_in(tile_1__5__11_cby_2__5__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__129_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_129_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__5__chanx_left_in(tile_1__6__11_sb_1__5__chanx_right_out[0:64]),
		.cby_2__6__chany_top_in(tile_1__2__129_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__6__13_ccff_tail),
		.sb_2__5__chanx_right_out(tile_2__6__11_sb_2__5__chanx_right_out[0:64]),
		.sb_2__5__chany_bottom_out(tile_2__6__11_sb_2__5__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_12__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__5__chanx_left_out(tile_2__6__11_cbx_2__5__chanx_left_out[0:64]),
		.cby_2__6__chany_top_out(tile_2__6__11_cby_2__6__chany_top_out[0:64]),
		.ccff_tail(tile_2__6__11_ccff_tail));

	tile_2__6_ tile_14__6_ (
		.prog_clk(prog_clk),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__14_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_2__5__chanx_right_in(tile_1__6__14_cbx_1__5__chanx_left_out[0:64]),
		.sb_2__5__chany_bottom_in(tile_1__5__12_cby_2__5__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__146_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_146_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__5__chanx_left_in(tile_1__6__12_sb_1__5__chanx_right_out[0:64]),
		.cby_2__6__chany_top_in(tile_1__2__146_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__6__12_ccff_tail),
		.sb_2__5__chanx_right_out(tile_2__6__12_sb_2__5__chanx_right_out[0:64]),
		.sb_2__5__chany_bottom_out(tile_2__6__12_sb_2__5__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_14__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__5__chanx_left_out(tile_2__6__12_cbx_2__5__chanx_left_out[0:64]),
		.cby_2__6__chany_top_out(tile_2__6__12_cby_2__6__chany_top_out[0:64]),
		.ccff_tail(tile_2__6__12_ccff_tail));

	tile_2__6_ tile_14__15_ (
		.prog_clk(prog_clk),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_1__5__15_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_2__5__chanx_right_in(tile_1__6__15_cbx_1__5__chanx_left_out[0:64]),
		.sb_2__5__chany_bottom_in(tile_1__5__13_cby_2__5__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__151_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_151_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__5__chanx_left_in(tile_1__6__13_sb_1__5__chanx_right_out[0:64]),
		.cby_2__6__chany_top_in(tile_1__2__151_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__6__15_ccff_tail),
		.sb_2__5__chanx_right_out(tile_2__6__13_sb_2__5__chanx_right_out[0:64]),
		.sb_2__5__chany_bottom_out(tile_2__6__13_sb_2__5__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_14__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__5__chanx_left_out(tile_2__6__13_cbx_2__5__chanx_left_out[0:64]),
		.cby_2__6__chany_top_out(tile_2__6__13_cby_2__6__chany_top_out[0:64]),
		.ccff_tail(tile_2__6__13_ccff_tail));

	tile_2__6_ tile_16__6_ (
		.prog_clk(prog_clk),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__16_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_2__5__chanx_right_in(tile_1__6__16_cbx_1__5__chanx_left_out[0:64]),
		.sb_2__5__chany_bottom_in(tile_1__5__14_cby_2__5__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__168_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_168_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__5__chanx_left_in(tile_1__6__14_sb_1__5__chanx_right_out[0:64]),
		.cby_2__6__chany_top_in(tile_1__2__168_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__6__14_ccff_tail),
		.sb_2__5__chanx_right_out(tile_2__6__14_sb_2__5__chanx_right_out[0:64]),
		.sb_2__5__chany_bottom_out(tile_2__6__14_sb_2__5__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__14_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__14_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_16__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__14_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__5__chanx_left_out(tile_2__6__14_cbx_2__5__chanx_left_out[0:64]),
		.cby_2__6__chany_top_out(tile_2__6__14_cby_2__6__chany_top_out[0:64]),
		.ccff_tail(tile_2__6__14_ccff_tail));

	tile_2__6_ tile_16__15_ (
		.prog_clk(prog_clk),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__6__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__6__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__6__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__6__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__6__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__5__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__6__17_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_2__5__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_2__5__chanx_right_in(tile_1__6__17_cbx_1__5__chanx_left_out[0:64]),
		.sb_2__5__chany_bottom_in(tile_1__5__15_cby_2__5__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__173_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_173_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__5__chanx_left_in(tile_1__6__15_sb_1__5__chanx_right_out[0:64]),
		.cby_2__6__chany_top_in(tile_1__2__173_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__6__17_ccff_tail),
		.sb_2__5__chanx_right_out(tile_2__6__15_sb_2__5__chanx_right_out[0:64]),
		.sb_2__5__chany_bottom_out(tile_2__6__15_sb_2__5__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__6__15_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__6__15_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_16__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__6__15_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__5__chanx_left_out(tile_2__6__15_cbx_2__5__chanx_left_out[0:64]),
		.cby_2__6__chany_top_out(tile_2__6__15_cby_2__6__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[24]));

	tile_2__11_ tile_2__11_ (
		.prog_clk(prog_clk),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__10__chanx_right_in(tile_1__11__1_cbx_1__10__chanx_left_out[0:64]),
		.sb_2__10__chany_bottom_in(tile_1__10__0_cby_2__10__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__17_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_17_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__10__chanx_left_in(tile_1__11__0_sb_1__10__chanx_right_out[0:64]),
		.cby_2__11__chany_top_in(tile_1__2__17_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__11__1_ccff_tail),
		.sb_2__10__chanx_right_out(tile_2__11__0_sb_2__10__chanx_right_out[0:64]),
		.sb_2__10__chany_bottom_out(tile_2__11__0_sb_2__10__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__11__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_2__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__11__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__10__chanx_left_out(tile_2__11__0_cbx_2__10__chanx_left_out[0:64]),
		.cby_2__11__chany_top_out(tile_2__11__0_cby_2__11__chany_top_out[0:64]),
		.ccff_tail(tile_2__11__0_ccff_tail));

	tile_2__11_ tile_4__11_ (
		.prog_clk(prog_clk),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__10__chanx_right_in(tile_1__11__2_cbx_1__10__chanx_left_out[0:64]),
		.sb_2__10__chany_bottom_in(tile_1__10__1_cby_2__10__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__39_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_39_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__10__chanx_left_in(tile_1__11__1_sb_1__10__chanx_right_out[0:64]),
		.cby_2__11__chany_top_in(tile_1__2__39_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__11__2_ccff_tail),
		.sb_2__10__chanx_right_out(tile_2__11__1_sb_2__10__chanx_right_out[0:64]),
		.sb_2__10__chany_bottom_out(tile_2__11__1_sb_2__10__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__11__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_4__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__11__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__10__chanx_left_out(tile_2__11__1_cbx_2__10__chanx_left_out[0:64]),
		.cby_2__11__chany_top_out(tile_2__11__1_cby_2__11__chany_top_out[0:64]),
		.ccff_tail(tile_2__11__1_ccff_tail));

	tile_2__11_ tile_6__11_ (
		.prog_clk(prog_clk),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__10__chanx_right_in(tile_1__11__3_cbx_1__10__chanx_left_out[0:64]),
		.sb_2__10__chany_bottom_in(tile_1__10__2_cby_2__10__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__61_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_61_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__10__chanx_left_in(tile_1__11__2_sb_1__10__chanx_right_out[0:64]),
		.cby_2__11__chany_top_in(tile_1__2__61_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__11__3_ccff_tail),
		.sb_2__10__chanx_right_out(tile_2__11__2_sb_2__10__chanx_right_out[0:64]),
		.sb_2__10__chany_bottom_out(tile_2__11__2_sb_2__10__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__11__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_6__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__11__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__10__chanx_left_out(tile_2__11__2_cbx_2__10__chanx_left_out[0:64]),
		.cby_2__11__chany_top_out(tile_2__11__2_cby_2__11__chany_top_out[0:64]),
		.ccff_tail(tile_2__11__2_ccff_tail));

	tile_2__11_ tile_8__11_ (
		.prog_clk(prog_clk),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__10__chanx_right_in(tile_1__11__4_cbx_1__10__chanx_left_out[0:64]),
		.sb_2__10__chany_bottom_in(tile_1__10__3_cby_2__10__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__83_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_83_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__10__chanx_left_in(tile_1__11__3_sb_1__10__chanx_right_out[0:64]),
		.cby_2__11__chany_top_in(tile_1__2__83_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__11__4_ccff_tail),
		.sb_2__10__chanx_right_out(tile_2__11__3_sb_2__10__chanx_right_out[0:64]),
		.sb_2__10__chany_bottom_out(tile_2__11__3_sb_2__10__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__11__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_8__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__11__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__10__chanx_left_out(tile_2__11__3_cbx_2__10__chanx_left_out[0:64]),
		.cby_2__11__chany_top_out(tile_2__11__3_cby_2__11__chany_top_out[0:64]),
		.ccff_tail(tile_2__11__3_ccff_tail));

	tile_2__11_ tile_10__11_ (
		.prog_clk(prog_clk),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__10__chanx_right_in(tile_1__11__5_cbx_1__10__chanx_left_out[0:64]),
		.sb_2__10__chany_bottom_in(tile_1__10__4_cby_2__10__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__105_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_105_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__10__chanx_left_in(tile_1__11__4_sb_1__10__chanx_right_out[0:64]),
		.cby_2__11__chany_top_in(tile_1__2__105_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[19]),
		.sb_2__10__chanx_right_out(tile_2__11__4_sb_2__10__chanx_right_out[0:64]),
		.sb_2__10__chany_bottom_out(tile_2__11__4_sb_2__10__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__11__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_10__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__11__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__10__chanx_left_out(tile_2__11__4_cbx_2__10__chanx_left_out[0:64]),
		.cby_2__11__chany_top_out(tile_2__11__4_cby_2__11__chany_top_out[0:64]),
		.ccff_tail(tile_2__11__4_ccff_tail));

	tile_2__11_ tile_12__11_ (
		.prog_clk(prog_clk),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__10__chanx_right_in(tile_1__11__6_cbx_1__10__chanx_left_out[0:64]),
		.sb_2__10__chany_bottom_in(tile_1__10__5_cby_2__10__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__127_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_127_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__10__chanx_left_in(tile_1__11__5_sb_1__10__chanx_right_out[0:64]),
		.cby_2__11__chany_top_in(tile_1__2__127_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__11__6_ccff_tail),
		.sb_2__10__chanx_right_out(tile_2__11__5_sb_2__10__chanx_right_out[0:64]),
		.sb_2__10__chany_bottom_out(tile_2__11__5_sb_2__10__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__11__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_12__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__11__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__10__chanx_left_out(tile_2__11__5_cbx_2__10__chanx_left_out[0:64]),
		.cby_2__11__chany_top_out(tile_2__11__5_cby_2__11__chany_top_out[0:64]),
		.ccff_tail(tile_2__11__5_ccff_tail));

	tile_2__11_ tile_14__11_ (
		.prog_clk(prog_clk),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__10__chanx_right_in(tile_1__11__7_cbx_1__10__chanx_left_out[0:64]),
		.sb_2__10__chany_bottom_in(tile_1__10__6_cby_2__10__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__149_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_149_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__10__chanx_left_in(tile_1__11__6_sb_1__10__chanx_right_out[0:64]),
		.cby_2__11__chany_top_in(tile_1__2__149_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__11__7_ccff_tail),
		.sb_2__10__chanx_right_out(tile_2__11__6_sb_2__10__chanx_right_out[0:64]),
		.sb_2__10__chany_bottom_out(tile_2__11__6_sb_2__10__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__11__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_14__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__11__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__10__chanx_left_out(tile_2__11__6_cbx_2__10__chanx_left_out[0:64]),
		.cby_2__11__chany_top_out(tile_2__11__6_cby_2__11__chany_top_out[0:64]),
		.ccff_tail(tile_2__11__6_ccff_tail));

	tile_2__11_ tile_16__11_ (
		.prog_clk(prog_clk),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__11__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__11__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__11__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__11__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__11__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_2__10__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__11__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_2__10__chanx_right_in(tile_1__11__8_cbx_1__10__chanx_left_out[0:64]),
		.sb_2__10__chany_bottom_in(tile_1__10__7_cby_2__10__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__171_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_171_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_2__10__chanx_left_in(tile_1__11__7_sb_1__10__chanx_right_out[0:64]),
		.cby_2__11__chany_top_in(tile_1__2__171_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__11__8_ccff_tail),
		.sb_2__10__chanx_right_out(tile_2__11__7_sb_2__10__chanx_right_out[0:64]),
		.sb_2__10__chany_bottom_out(tile_2__11__7_sb_2__10__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_2__11__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_2__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_2__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_2__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_2__11__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_16__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_2__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_2__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_2__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_2__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_2__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_2__11__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_2__10__chanx_left_out(tile_2__11__7_cbx_2__10__chanx_left_out[0:64]),
		.cby_2__11__chany_top_out(tile_2__11__7_cby_2__11__chany_top_out[0:64]),
		.ccff_tail(tile_2__11__7_ccff_tail));

	tile_17__5_ tile_17__5_ (
		.prog_clk(prog_clk),
		.sb_17__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_17__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_17__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_17__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_17__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_17__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_17__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__178_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_17__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__178_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_17__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__178_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_17__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__178_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_17__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_17__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_17__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_17__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_17__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_17__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__178_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_18__4__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__13_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__4__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__13_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__4__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__14_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__4__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__14_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_18__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_18__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_18__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_18__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_18__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_18__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_18__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_18__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_18__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_17__4__chany_bottom_in(tile_1__2__178_cby_1__2__chany_top_out[0:64]),
		.sb_18__4__chany_bottom_in(tile_18__2__2_cby_18__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__16_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_17__4__chanx_left_in(tile_1__5__14_sb_2__4__chanx_right_out[0:64]),
		.cby_18__5__chany_top_in(tile_18__6__0_sb_18__5__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[9]),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_17__5__0_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cby_18__5__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_17__5__0_cby_18__5__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_18__5__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_17__5__0_cby_18__5__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_17__4__chany_bottom_out(tile_17__5__0_sb_17__4__chany_bottom_out[0:64]),
		.sb_18__4__chany_bottom_out(tile_17__5__0_sb_18__4__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_17__5__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_17__4__chanx_left_out(tile_17__5__0_cbx_17__4__chanx_left_out[0:64]),
		.cby_18__5__chany_top_out(tile_17__5__0_cby_18__5__chany_top_out[0:64]),
		.ccff_tail(tile_17__5__0_ccff_tail));

	tile_17__5_ tile_17__14_ (
		.prog_clk(prog_clk),
		.sb_17__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_17__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_17__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_17__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_17__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_17__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_17__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__183_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_17__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__183_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_17__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__183_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_17__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__183_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_17__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_17__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_17__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_17__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_17__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_17__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__183_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_18__4__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__4_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__4__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__4_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__4__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__5_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__4__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__5_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_18__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_18__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_18__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_18__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_18__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_18__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_18__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_18__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_18__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_17__4__chany_bottom_in(tile_1__2__183_cby_1__2__chany_top_out[0:64]),
		.sb_18__4__chany_bottom_in(tile_18__2__7_cby_18__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_1__6__17_cbx_1__5__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_17__4__chanx_left_in(tile_1__5__15_sb_2__4__chanx_right_out[0:64]),
		.cby_18__5__chany_top_in(tile_18__6__2_sb_18__5__chany_bottom_out[0:64]),
		.ccff_head(tile_1__5__15_ccff_tail),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_17__5__1_cbx_17__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cby_18__5__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_17__5__1_cby_18__5__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_18__5__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_17__5__1_cby_18__5__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_17__4__chany_bottom_out(tile_17__5__1_sb_17__4__chany_bottom_out[0:64]),
		.sb_18__4__chany_bottom_out(tile_17__5__1_sb_18__4__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_17__5__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_17__4__chanx_left_out(tile_17__5__1_cbx_17__4__chanx_left_out[0:64]),
		.cby_18__5__chany_top_out(tile_17__5__1_cby_18__5__chany_top_out[0:64]),
		.ccff_tail(tile_17__5__1_ccff_tail));

	tile_17__10_ tile_17__10_ (
		.prog_clk(prog_clk),
		.sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_17__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__181_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_17__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__181_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_17__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__181_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_17__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__181_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__181_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_18__9__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__8_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__9__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__8_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__9__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__9_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__9__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__9_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_18__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_18__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_18__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_17__9__chany_bottom_in(tile_1__2__181_cby_1__2__chany_top_out[0:64]),
		.sb_18__9__chany_bottom_in(tile_18__2__5_cby_18__2__chany_top_out[0:64]),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_(tile_1__11__8_cbx_1__10__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.cbx_17__9__chanx_left_in(tile_1__10__7_sb_2__9__chanx_right_out[0:64]),
		.cby_18__10__chany_top_in(tile_18__6__1_sb_18__5__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[18]),
		.cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_17__10__0_cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cby_18__10__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_17__10__0_cby_18__10__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_18__10__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_17__10__0_cby_18__10__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_17__9__chany_bottom_out(tile_17__10__0_sb_17__9__chany_bottom_out[0:64]),
		.sb_18__9__chany_bottom_out(tile_17__10__0_sb_18__9__chany_bottom_out[0:64]),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_17__10__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.cbx_17__9__chanx_left_out(tile_17__10__0_cbx_17__9__chanx_left_out[0:64]),
		.cby_18__10__chany_top_out(tile_17__10__0_cby_18__10__chany_top_out[0:64]),
		.ccff_tail(tile_17__10__0_ccff_tail));

	tile_18__1_ tile_18__1_ (
		.prog_clk(prog_clk),
		.sb_18__0__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__17_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__0__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__17_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__0_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__0_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_187_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_18__0__chanx_left_in(tile_1__1__16_sb_1__0__chanx_right_out[0:64]),
		.cby_18__1__chany_top_in(tile_18__2__0_sb_18__1__chany_bottom_out[0:64]),
		.ccff_head(tile_19__1__17_ccff_tail),
		.cbx_18__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__1__0_cbx_18__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_18__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__1__0_cbx_18__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.cby_18__1__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__1__0_cby_18__1__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_18__1__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__1__0_cby_18__1__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_18__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_18__0__chanx_left_out(tile_18__1__0_cbx_18__0__chanx_left_out[0:64]),
		.cby_18__1__chany_top_out(tile_18__1__0_cby_18__1__chany_top_out[0:64]),
		.ccff_tail(tile_18__1__0_ccff_tail));

	tile_18__2_ tile_18__2_ (
		.prog_clk(prog_clk),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__16_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__16_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__17_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__17_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_18__1__chany_bottom_in(tile_18__1__0_cby_18__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_188_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_18__1__chanx_left_in(tile_1__2__176_sb_1__1__chanx_right_out[0:64]),
		.cby_18__2__chany_top_in(tile_18__2__1_sb_18__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__176_ccff_tail),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__0_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__0_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__0_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_18__1__chany_bottom_out(tile_18__2__0_sb_18__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_18__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_18__1__chanx_left_out(tile_18__2__0_cbx_18__1__chanx_left_out[0:64]),
		.cby_18__2__chany_top_out(tile_18__2__0_cby_18__2__chany_top_out[0:64]),
		.ccff_tail(tile_18__2__0_ccff_tail));

	tile_18__2_ tile_18__3_ (
		.prog_clk(prog_clk),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__15_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__15_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__16_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__16_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_18__1__chany_bottom_in(tile_18__2__0_cby_18__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_189_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_18__1__chanx_left_in(tile_1__2__177_sb_1__1__chanx_right_out[0:64]),
		.cby_18__2__chany_top_in(tile_18__2__2_sb_18__1__chany_bottom_out[0:64]),
		.ccff_head(tile_19__1__15_ccff_tail),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__1_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__1_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__1_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_18__1__chany_bottom_out(tile_18__2__1_sb_18__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_18__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_18__1__chanx_left_out(tile_18__2__1_cbx_18__1__chanx_left_out[0:64]),
		.cby_18__2__chany_top_out(tile_18__2__1_cby_18__2__chany_top_out[0:64]),
		.ccff_tail(tile_18__2__1_ccff_tail));

	tile_18__2_ tile_18__4_ (
		.prog_clk(prog_clk),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__14_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__14_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__15_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__15_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_18__1__chany_bottom_in(tile_18__2__1_cby_18__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_17__5__0_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_18__4__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_18__1__chanx_left_in(tile_1__2__178_sb_1__1__chanx_right_out[0:64]),
		.cby_18__2__chany_top_in(tile_17__5__0_sb_18__4__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__178_ccff_tail),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__2_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__2_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__2_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_18__1__chany_bottom_out(tile_18__2__2_sb_18__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_18__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_18__1__chanx_left_out(tile_18__2__2_cbx_18__1__chanx_left_out[0:64]),
		.cby_18__2__chany_top_out(tile_18__2__2_cby_18__2__chany_top_out[0:64]),
		.ccff_tail(tile_18__2__2_ccff_tail));

	tile_18__2_ tile_18__7_ (
		.prog_clk(prog_clk),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__11_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__11_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__12_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__12_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_18__1__chany_bottom_in(tile_18__6__0_cby_18__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_191_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_18__1__chanx_left_in(tile_1__2__179_sb_1__1__chanx_right_out[0:64]),
		.cby_18__2__chany_top_in(tile_18__2__4_sb_18__1__chany_bottom_out[0:64]),
		.ccff_head(tile_19__1__11_ccff_tail),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__3_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__3_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_18__1__chany_bottom_out(tile_18__2__3_sb_18__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_18__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_18__1__chanx_left_out(tile_18__2__3_cbx_18__1__chanx_left_out[0:64]),
		.cby_18__2__chany_top_out(tile_18__2__3_cby_18__2__chany_top_out[0:64]),
		.ccff_tail(tile_18__2__3_ccff_tail));

	tile_18__2_ tile_18__8_ (
		.prog_clk(prog_clk),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__10_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__10_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__11_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__11_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_18__1__chany_bottom_in(tile_18__2__3_cby_18__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_192_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_18__1__chanx_left_in(tile_1__2__180_sb_1__1__chanx_right_out[0:64]),
		.cby_18__2__chany_top_in(tile_18__2__5_sb_18__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__180_ccff_tail),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__4_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__4_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__4_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_18__1__chany_bottom_out(tile_18__2__4_sb_18__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_18__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_18__1__chanx_left_out(tile_18__2__4_cbx_18__1__chanx_left_out[0:64]),
		.cby_18__2__chany_top_out(tile_18__2__4_cby_18__2__chany_top_out[0:64]),
		.ccff_tail(tile_18__2__4_ccff_tail));

	tile_18__2_ tile_18__9_ (
		.prog_clk(prog_clk),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__9_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__9_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__10_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__10_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_18__1__chany_bottom_in(tile_18__2__4_cby_18__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_17__10__0_cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_18__9__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_18__1__chanx_left_in(tile_1__2__181_sb_1__1__chanx_right_out[0:64]),
		.cby_18__2__chany_top_in(tile_17__10__0_sb_18__9__chany_bottom_out[0:64]),
		.ccff_head(tile_19__1__9_ccff_tail),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__5_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__5_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__5_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_18__1__chany_bottom_out(tile_18__2__5_sb_18__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_18__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_18__1__chanx_left_out(tile_18__2__5_cbx_18__1__chanx_left_out[0:64]),
		.cby_18__2__chany_top_out(tile_18__2__5_cby_18__2__chany_top_out[0:64]),
		.ccff_tail(tile_18__2__5_ccff_tail));

	tile_18__2_ tile_18__12_ (
		.prog_clk(prog_clk),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__6_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__6_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__7_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__7_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_18__1__chany_bottom_in(tile_18__6__1_cby_18__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_194_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_18__1__chanx_left_in(tile_1__2__182_sb_1__1__chanx_right_out[0:64]),
		.cby_18__2__chany_top_in(tile_18__2__7_sb_18__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__182_ccff_tail),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__6_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__6_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_18__1__chany_bottom_out(tile_18__2__6_sb_18__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_18__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_18__1__chanx_left_out(tile_18__2__6_cbx_18__1__chanx_left_out[0:64]),
		.cby_18__2__chany_top_out(tile_18__2__6_cby_18__2__chany_top_out[0:64]),
		.ccff_tail(tile_18__2__6_ccff_tail));

	tile_18__2_ tile_18__13_ (
		.prog_clk(prog_clk),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__5_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__5_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__6_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__6_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_18__1__chany_bottom_in(tile_18__2__6_cby_18__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_17__5__1_cbx_18__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_18__13__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_18__1__chanx_left_in(tile_1__2__183_sb_1__1__chanx_right_out[0:64]),
		.cby_18__2__chany_top_in(tile_17__5__1_sb_18__4__chany_bottom_out[0:64]),
		.ccff_head(tile_19__1__5_ccff_tail),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__7_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__7_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__7_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_18__1__chany_bottom_out(tile_18__2__7_sb_18__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_18__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_18__1__chanx_left_out(tile_18__2__7_cbx_18__1__chanx_left_out[0:64]),
		.cby_18__2__chany_top_out(tile_18__2__7_cby_18__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[21]));

	tile_18__2_ tile_18__16_ (
		.prog_clk(prog_clk),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__2_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__2_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__3_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__3_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_18__1__chany_bottom_in(tile_18__6__2_cby_18__6__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_196_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_18__1__chanx_left_in(tile_1__2__184_sb_1__1__chanx_right_out[0:64]),
		.cby_18__2__chany_top_in(tile_18__2__9_sb_18__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__184_ccff_tail),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__8_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__8_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_18__1__chany_bottom_out(tile_18__2__8_sb_18__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_18__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_18__1__chanx_left_out(tile_18__2__8_cbx_18__1__chanx_left_out[0:64]),
		.cby_18__2__chany_top_out(tile_18__2__8_cby_18__2__chany_top_out[0:64]),
		.ccff_tail(tile_18__2__8_ccff_tail));

	tile_18__2_ tile_18__17_ (
		.prog_clk(prog_clk),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__1_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__1_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__2_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__2_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_18__1__chany_bottom_in(tile_18__2__8_cby_18__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_197_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_18__1__chanx_left_in(tile_1__2__185_sb_1__1__chanx_right_out[0:64]),
		.cby_18__2__chany_top_in(tile_18__2__10_sb_18__1__chany_bottom_out[0:64]),
		.ccff_head(tile_19__1__1_ccff_tail),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__9_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__9_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__9_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_18__1__chany_bottom_out(tile_18__2__9_sb_18__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_18__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_18__1__chanx_left_out(tile_18__2__9_cbx_18__1__chanx_left_out[0:64]),
		.cby_18__2__chany_top_out(tile_18__2__9_cby_18__2__chany_top_out[0:64]),
		.ccff_tail(tile_18__2__9_ccff_tail));

	tile_18__2_ tile_18__18_ (
		.prog_clk(prog_clk),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__0_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__0_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__1_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__1__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__1_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_18__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_18__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_18__1__chany_bottom_in(tile_18__2__9_cby_18__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__19__0_cbx_18__18__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_18__18__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_18__1__chanx_left_in(tile_1__2__186_sb_1__1__chanx_right_out[0:64]),
		.cby_18__2__chany_top_in(tile_18__19__0_sb_18__18__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__186_ccff_tail),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__10_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__2__10_cby_18__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__2__10_cby_18__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_18__1__chany_bottom_out(tile_18__2__10_sb_18__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_18__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_18__1__chanx_left_out(tile_18__2__10_cbx_18__1__chanx_left_out[0:64]),
		.cby_18__2__chany_top_out(tile_18__2__10_cby_18__2__chany_top_out[0:64]),
		.ccff_tail(tile_18__2__10_ccff_tail));

	tile_18__6_ tile_18__6_ (
		.prog_clk(prog_clk),
		.sb_18__5__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__12_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__5__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__12_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__5__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__13_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__5__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__13_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__5__chany_bottom_in(tile_17__5__0_cby_18__5__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__3_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_190_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_18__5__chanx_left_in(tile_1__6__16_sb_1__5__chanx_right_out[0:64]),
		.cby_18__6__chany_top_in(tile_18__2__3_sb_18__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__6__16_ccff_tail),
		.cby_18__6__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__6__0_cby_18__6__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_18__6__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__6__0_cby_18__6__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_18__5__chany_bottom_out(tile_18__6__0_sb_18__5__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__6__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__6__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_18__6__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__6__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_18__5__chanx_left_out(tile_18__6__0_cbx_18__5__chanx_left_out[0:64]),
		.cby_18__6__chany_top_out(tile_18__6__0_cby_18__6__chany_top_out[0:64]),
		.ccff_tail(tile_18__6__0_ccff_tail));

	tile_18__6_ tile_18__11_ (
		.prog_clk(prog_clk),
		.sb_18__5__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__7_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__5__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__7_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__5__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__8_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__5__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__8_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__5__chany_bottom_in(tile_17__10__0_cby_18__10__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__6_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_193_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_18__5__chanx_left_in(tile_1__11__8_sb_1__10__chanx_right_out[0:64]),
		.cby_18__6__chany_top_in(tile_18__2__6_sb_18__1__chany_bottom_out[0:64]),
		.ccff_head(tile_19__1__7_ccff_tail),
		.cby_18__6__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__6__1_cby_18__6__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_18__6__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__6__1_cby_18__6__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_18__5__chany_bottom_out(tile_18__6__1_sb_18__5__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__6__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__6__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_18__11__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__6__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_18__5__chanx_left_out(tile_18__6__1_cbx_18__5__chanx_left_out[0:64]),
		.cby_18__6__chany_top_out(tile_18__6__1_cby_18__6__chany_top_out[0:64]),
		.ccff_tail(tile_18__6__1_ccff_tail));

	tile_18__6_ tile_18__15_ (
		.prog_clk(prog_clk),
		.sb_18__5__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__3_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__5__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__3_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__5__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_19__1__4_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_18__5__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_19__1__4_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_18__5__chany_bottom_in(tile_17__5__1_cby_18__5__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_18__2__8_cbx_18__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_195_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk_i),
		.cbx_18__5__chanx_left_in(tile_1__6__17_sb_1__5__chanx_right_out[0:64]),
		.cby_18__6__chany_top_in(tile_18__2__8_sb_18__1__chany_bottom_out[0:64]),
		.ccff_head(tile_19__1__3_ccff_tail),
		.cby_18__6__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_18__6__2_cby_18__6__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_18__6__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_18__6__2_cby_18__6__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_18__5__chany_bottom_out(tile_18__6__2_sb_18__5__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_18__6__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_18__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_18__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_18__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_18__6__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_18__15__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_18__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_18__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_18__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_18__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_18__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_18__6__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_18__5__chanx_left_out(tile_18__6__2_cbx_18__5__chanx_left_out[0:64]),
		.cby_18__6__chany_top_out(tile_18__6__2_cby_18__6__chany_top_out[0:64]),
		.ccff_tail(tile_18__6__2_ccff_tail));

	direct_interc direct_interc_0_ (
		.in(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_0_out));

	direct_interc direct_interc_1_ (
		.in(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_1_out));

	direct_interc direct_interc_2_ (
		.in(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_2_out));

	direct_interc direct_interc_3_ (
		.in(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_3_out));

	direct_interc direct_interc_4_ (
		.in(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_4_out));

	direct_interc direct_interc_5_ (
		.in(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_5_out));

	direct_interc direct_interc_6_ (
		.in(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_6_out));

	direct_interc direct_interc_7_ (
		.in(tile_1__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_7_out));

	direct_interc direct_interc_8_ (
		.in(tile_1__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_8_out));

	direct_interc direct_interc_9_ (
		.in(tile_1__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_9_out));

	direct_interc direct_interc_10_ (
		.in(tile_1__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_10_out));

	direct_interc direct_interc_11_ (
		.in(tile_1__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_11_out));

	direct_interc direct_interc_12_ (
		.in(tile_1__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_12_out));

	direct_interc direct_interc_13_ (
		.in(tile_1__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_13_out));

	direct_interc direct_interc_14_ (
		.in(tile_1__2__14_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_14_out));

	direct_interc direct_interc_15_ (
		.in(tile_1__2__15_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_15_out));

	direct_interc direct_interc_16_ (
		.in(tile_1__2__16_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_16_out));

	direct_interc direct_interc_17_ (
		.in(tile_1__2__17_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_17_out));

	direct_interc direct_interc_18_ (
		.in(tile_1__2__18_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_18_out));

	direct_interc direct_interc_19_ (
		.in(tile_1__2__19_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_19_out));

	direct_interc direct_interc_20_ (
		.in(tile_1__2__20_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_20_out));

	direct_interc direct_interc_21_ (
		.in(tile_1__2__21_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_21_out));

	direct_interc direct_interc_22_ (
		.in(tile_1__2__22_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_22_out));

	direct_interc direct_interc_23_ (
		.in(tile_1__2__23_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_23_out));

	direct_interc direct_interc_24_ (
		.in(tile_1__2__24_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_24_out));

	direct_interc direct_interc_25_ (
		.in(tile_1__2__25_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_25_out));

	direct_interc direct_interc_26_ (
		.in(tile_1__2__26_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_26_out));

	direct_interc direct_interc_27_ (
		.in(tile_1__2__27_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_27_out));

	direct_interc direct_interc_28_ (
		.in(tile_1__2__28_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_28_out));

	direct_interc direct_interc_29_ (
		.in(tile_1__2__29_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_29_out));

	direct_interc direct_interc_30_ (
		.in(tile_1__2__30_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_30_out));

	direct_interc direct_interc_31_ (
		.in(tile_1__2__31_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_31_out));

	direct_interc direct_interc_32_ (
		.in(tile_1__2__32_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_32_out));

	direct_interc direct_interc_33_ (
		.in(tile_1__2__33_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_33_out));

	direct_interc direct_interc_34_ (
		.in(tile_1__2__34_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_34_out));

	direct_interc direct_interc_35_ (
		.in(tile_1__2__35_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_35_out));

	direct_interc direct_interc_36_ (
		.in(tile_1__2__36_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_36_out));

	direct_interc direct_interc_37_ (
		.in(tile_1__2__37_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_37_out));

	direct_interc direct_interc_38_ (
		.in(tile_1__2__38_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_38_out));

	direct_interc direct_interc_39_ (
		.in(tile_1__2__39_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_39_out));

	direct_interc direct_interc_40_ (
		.in(tile_1__2__40_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_40_out));

	direct_interc direct_interc_41_ (
		.in(tile_1__2__41_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_41_out));

	direct_interc direct_interc_42_ (
		.in(tile_1__2__42_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_42_out));

	direct_interc direct_interc_43_ (
		.in(tile_1__2__43_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_43_out));

	direct_interc direct_interc_44_ (
		.in(tile_1__2__44_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_44_out));

	direct_interc direct_interc_45_ (
		.in(tile_1__2__45_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_45_out));

	direct_interc direct_interc_46_ (
		.in(tile_1__2__46_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_46_out));

	direct_interc direct_interc_47_ (
		.in(tile_1__2__47_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_47_out));

	direct_interc direct_interc_48_ (
		.in(tile_1__2__48_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_48_out));

	direct_interc direct_interc_49_ (
		.in(tile_1__2__49_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_49_out));

	direct_interc direct_interc_50_ (
		.in(tile_1__2__50_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_50_out));

	direct_interc direct_interc_51_ (
		.in(tile_1__2__51_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_51_out));

	direct_interc direct_interc_52_ (
		.in(tile_1__2__52_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_52_out));

	direct_interc direct_interc_53_ (
		.in(tile_1__2__53_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_53_out));

	direct_interc direct_interc_54_ (
		.in(tile_1__2__54_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_54_out));

	direct_interc direct_interc_55_ (
		.in(tile_1__2__55_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_55_out));

	direct_interc direct_interc_56_ (
		.in(tile_1__2__56_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_56_out));

	direct_interc direct_interc_57_ (
		.in(tile_1__2__57_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_57_out));

	direct_interc direct_interc_58_ (
		.in(tile_1__2__58_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_58_out));

	direct_interc direct_interc_59_ (
		.in(tile_1__2__59_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_59_out));

	direct_interc direct_interc_60_ (
		.in(tile_1__2__60_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_60_out));

	direct_interc direct_interc_61_ (
		.in(tile_1__2__61_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_61_out));

	direct_interc direct_interc_62_ (
		.in(tile_1__2__62_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_62_out));

	direct_interc direct_interc_63_ (
		.in(tile_1__2__63_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_63_out));

	direct_interc direct_interc_64_ (
		.in(tile_1__2__64_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_64_out));

	direct_interc direct_interc_65_ (
		.in(tile_1__2__65_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_65_out));

	direct_interc direct_interc_66_ (
		.in(tile_1__2__66_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_66_out));

	direct_interc direct_interc_67_ (
		.in(tile_1__2__67_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_67_out));

	direct_interc direct_interc_68_ (
		.in(tile_1__2__68_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_68_out));

	direct_interc direct_interc_69_ (
		.in(tile_1__2__69_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_69_out));

	direct_interc direct_interc_70_ (
		.in(tile_1__2__70_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_70_out));

	direct_interc direct_interc_71_ (
		.in(tile_1__2__71_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_71_out));

	direct_interc direct_interc_72_ (
		.in(tile_1__2__72_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_72_out));

	direct_interc direct_interc_73_ (
		.in(tile_1__2__73_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_73_out));

	direct_interc direct_interc_74_ (
		.in(tile_1__2__74_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_74_out));

	direct_interc direct_interc_75_ (
		.in(tile_1__2__75_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_75_out));

	direct_interc direct_interc_76_ (
		.in(tile_1__2__76_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_76_out));

	direct_interc direct_interc_77_ (
		.in(tile_1__2__77_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_77_out));

	direct_interc direct_interc_78_ (
		.in(tile_1__2__78_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_78_out));

	direct_interc direct_interc_79_ (
		.in(tile_1__2__79_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_79_out));

	direct_interc direct_interc_80_ (
		.in(tile_1__2__80_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_80_out));

	direct_interc direct_interc_81_ (
		.in(tile_1__2__81_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_81_out));

	direct_interc direct_interc_82_ (
		.in(tile_1__2__82_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_82_out));

	direct_interc direct_interc_83_ (
		.in(tile_1__2__83_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_83_out));

	direct_interc direct_interc_84_ (
		.in(tile_1__2__84_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_84_out));

	direct_interc direct_interc_85_ (
		.in(tile_1__2__85_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_85_out));

	direct_interc direct_interc_86_ (
		.in(tile_1__2__86_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_86_out));

	direct_interc direct_interc_87_ (
		.in(tile_1__2__87_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_87_out));

	direct_interc direct_interc_88_ (
		.in(tile_1__2__88_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_88_out));

	direct_interc direct_interc_89_ (
		.in(tile_1__2__89_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_89_out));

	direct_interc direct_interc_90_ (
		.in(tile_1__2__90_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_90_out));

	direct_interc direct_interc_91_ (
		.in(tile_1__2__91_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_91_out));

	direct_interc direct_interc_92_ (
		.in(tile_1__2__92_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_92_out));

	direct_interc direct_interc_93_ (
		.in(tile_1__2__93_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_93_out));

	direct_interc direct_interc_94_ (
		.in(tile_1__2__94_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_94_out));

	direct_interc direct_interc_95_ (
		.in(tile_1__2__95_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_95_out));

	direct_interc direct_interc_96_ (
		.in(tile_1__2__96_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_96_out));

	direct_interc direct_interc_97_ (
		.in(tile_1__2__97_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_97_out));

	direct_interc direct_interc_98_ (
		.in(tile_1__2__98_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_98_out));

	direct_interc direct_interc_99_ (
		.in(tile_1__2__99_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_99_out));

	direct_interc direct_interc_100_ (
		.in(tile_1__2__100_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_100_out));

	direct_interc direct_interc_101_ (
		.in(tile_1__2__101_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_101_out));

	direct_interc direct_interc_102_ (
		.in(tile_1__2__102_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_102_out));

	direct_interc direct_interc_103_ (
		.in(tile_1__2__103_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_103_out));

	direct_interc direct_interc_104_ (
		.in(tile_1__2__104_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_104_out));

	direct_interc direct_interc_105_ (
		.in(tile_1__2__105_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_105_out));

	direct_interc direct_interc_106_ (
		.in(tile_1__2__106_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_106_out));

	direct_interc direct_interc_107_ (
		.in(tile_1__2__107_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_107_out));

	direct_interc direct_interc_108_ (
		.in(tile_1__2__108_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_108_out));

	direct_interc direct_interc_109_ (
		.in(tile_1__2__109_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_109_out));

	direct_interc direct_interc_110_ (
		.in(tile_1__2__110_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_110_out));

	direct_interc direct_interc_111_ (
		.in(tile_1__2__111_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_111_out));

	direct_interc direct_interc_112_ (
		.in(tile_1__2__112_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_112_out));

	direct_interc direct_interc_113_ (
		.in(tile_1__2__113_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_113_out));

	direct_interc direct_interc_114_ (
		.in(tile_1__2__114_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_114_out));

	direct_interc direct_interc_115_ (
		.in(tile_1__2__115_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_115_out));

	direct_interc direct_interc_116_ (
		.in(tile_1__2__116_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_116_out));

	direct_interc direct_interc_117_ (
		.in(tile_1__2__117_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_117_out));

	direct_interc direct_interc_118_ (
		.in(tile_1__2__118_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_118_out));

	direct_interc direct_interc_119_ (
		.in(tile_1__2__119_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_119_out));

	direct_interc direct_interc_120_ (
		.in(tile_1__2__120_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_120_out));

	direct_interc direct_interc_121_ (
		.in(tile_1__2__121_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_121_out));

	direct_interc direct_interc_122_ (
		.in(tile_1__2__122_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_122_out));

	direct_interc direct_interc_123_ (
		.in(tile_1__2__123_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_123_out));

	direct_interc direct_interc_124_ (
		.in(tile_1__2__124_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_124_out));

	direct_interc direct_interc_125_ (
		.in(tile_1__2__125_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_125_out));

	direct_interc direct_interc_126_ (
		.in(tile_1__2__126_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_126_out));

	direct_interc direct_interc_127_ (
		.in(tile_1__2__127_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_127_out));

	direct_interc direct_interc_128_ (
		.in(tile_1__2__128_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_128_out));

	direct_interc direct_interc_129_ (
		.in(tile_1__2__129_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_129_out));

	direct_interc direct_interc_130_ (
		.in(tile_1__2__130_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_130_out));

	direct_interc direct_interc_131_ (
		.in(tile_1__2__131_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_131_out));

	direct_interc direct_interc_132_ (
		.in(tile_1__2__132_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_132_out));

	direct_interc direct_interc_133_ (
		.in(tile_1__2__133_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_133_out));

	direct_interc direct_interc_134_ (
		.in(tile_1__2__134_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_134_out));

	direct_interc direct_interc_135_ (
		.in(tile_1__2__135_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_135_out));

	direct_interc direct_interc_136_ (
		.in(tile_1__2__136_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_136_out));

	direct_interc direct_interc_137_ (
		.in(tile_1__2__137_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_137_out));

	direct_interc direct_interc_138_ (
		.in(tile_1__2__138_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_138_out));

	direct_interc direct_interc_139_ (
		.in(tile_1__2__139_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_139_out));

	direct_interc direct_interc_140_ (
		.in(tile_1__2__140_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_140_out));

	direct_interc direct_interc_141_ (
		.in(tile_1__2__141_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_141_out));

	direct_interc direct_interc_142_ (
		.in(tile_1__2__142_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_142_out));

	direct_interc direct_interc_143_ (
		.in(tile_1__2__143_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_143_out));

	direct_interc direct_interc_144_ (
		.in(tile_1__2__144_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_144_out));

	direct_interc direct_interc_145_ (
		.in(tile_1__2__145_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_145_out));

	direct_interc direct_interc_146_ (
		.in(tile_1__2__146_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_146_out));

	direct_interc direct_interc_147_ (
		.in(tile_1__2__147_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_147_out));

	direct_interc direct_interc_148_ (
		.in(tile_1__2__148_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_148_out));

	direct_interc direct_interc_149_ (
		.in(tile_1__2__149_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_149_out));

	direct_interc direct_interc_150_ (
		.in(tile_1__2__150_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_150_out));

	direct_interc direct_interc_151_ (
		.in(tile_1__2__151_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_151_out));

	direct_interc direct_interc_152_ (
		.in(tile_1__2__152_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_152_out));

	direct_interc direct_interc_153_ (
		.in(tile_1__2__153_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_153_out));

	direct_interc direct_interc_154_ (
		.in(tile_1__2__154_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_154_out));

	direct_interc direct_interc_155_ (
		.in(tile_1__2__155_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_155_out));

	direct_interc direct_interc_156_ (
		.in(tile_1__2__156_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_156_out));

	direct_interc direct_interc_157_ (
		.in(tile_1__2__157_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_157_out));

	direct_interc direct_interc_158_ (
		.in(tile_1__2__158_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_158_out));

	direct_interc direct_interc_159_ (
		.in(tile_1__2__159_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_159_out));

	direct_interc direct_interc_160_ (
		.in(tile_1__2__160_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_160_out));

	direct_interc direct_interc_161_ (
		.in(tile_1__2__161_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_161_out));

	direct_interc direct_interc_162_ (
		.in(tile_1__2__162_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_162_out));

	direct_interc direct_interc_163_ (
		.in(tile_1__2__163_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_163_out));

	direct_interc direct_interc_164_ (
		.in(tile_1__2__164_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_164_out));

	direct_interc direct_interc_165_ (
		.in(tile_1__2__165_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_165_out));

	direct_interc direct_interc_166_ (
		.in(tile_1__2__166_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_166_out));

	direct_interc direct_interc_167_ (
		.in(tile_1__2__167_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_167_out));

	direct_interc direct_interc_168_ (
		.in(tile_1__2__168_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_168_out));

	direct_interc direct_interc_169_ (
		.in(tile_1__2__169_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_169_out));

	direct_interc direct_interc_170_ (
		.in(tile_1__2__170_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_170_out));

	direct_interc direct_interc_171_ (
		.in(tile_1__2__171_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_171_out));

	direct_interc direct_interc_172_ (
		.in(tile_1__2__172_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_172_out));

	direct_interc direct_interc_173_ (
		.in(tile_1__2__173_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_173_out));

	direct_interc direct_interc_174_ (
		.in(tile_1__2__174_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_174_out));

	direct_interc direct_interc_175_ (
		.in(tile_1__2__175_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_175_out));

	direct_interc direct_interc_176_ (
		.in(tile_1__2__176_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_176_out));

	direct_interc direct_interc_177_ (
		.in(tile_1__2__177_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_177_out));

	direct_interc direct_interc_178_ (
		.in(tile_1__2__178_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_178_out));

	direct_interc direct_interc_179_ (
		.in(tile_1__2__179_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_179_out));

	direct_interc direct_interc_180_ (
		.in(tile_1__2__180_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_180_out));

	direct_interc direct_interc_181_ (
		.in(tile_1__2__181_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_181_out));

	direct_interc direct_interc_182_ (
		.in(tile_1__2__182_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_182_out));

	direct_interc direct_interc_183_ (
		.in(tile_1__2__183_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_183_out));

	direct_interc direct_interc_184_ (
		.in(tile_1__2__184_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_184_out));

	direct_interc direct_interc_185_ (
		.in(tile_1__2__185_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_185_out));

	direct_interc direct_interc_186_ (
		.in(tile_1__2__186_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_186_out));

	direct_interc direct_interc_187_ (
		.in(tile_18__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_187_out));

	direct_interc direct_interc_188_ (
		.in(tile_18__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_188_out));

	direct_interc direct_interc_189_ (
		.in(tile_18__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_189_out));

	direct_interc direct_interc_190_ (
		.in(tile_18__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_190_out));

	direct_interc direct_interc_191_ (
		.in(tile_18__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_191_out));

	direct_interc direct_interc_192_ (
		.in(tile_18__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_192_out));

	direct_interc direct_interc_193_ (
		.in(tile_18__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_193_out));

	direct_interc direct_interc_194_ (
		.in(tile_18__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_194_out));

	direct_interc direct_interc_195_ (
		.in(tile_18__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_195_out));

	direct_interc direct_interc_196_ (
		.in(tile_18__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_196_out));

	direct_interc direct_interc_197_ (
		.in(tile_18__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_197_out));

endmodule
// ----- END Verilog module for fpga_top -----

//----- Default net type -----
`default_nettype wire




