/*verilator tracing_off*/
//Example
//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[1][4]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed Aug 14 09:11:36 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype wire

// ----- Verilog module for sb_1__4_ -----
module sb_1__4_(prog_clk,
                chanx_right_in,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_,
                chany_bottom_in,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_,
                chanx_left_in,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_,
                ccff_head,
                chanx_right_out,
                chany_bottom_out,
                chanx_left_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:64] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_;
//----- INPUT PORTS -----
input [0:64] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
//----- INPUT PORTS -----
input [0:64] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:64] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:64] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:64] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_tree_tapbuf_size2_0_sram;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_10_sram;
wire [0:1] mux_tree_tapbuf_size2_10_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_11_sram;
wire [0:1] mux_tree_tapbuf_size2_11_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_12_sram;
wire [0:1] mux_tree_tapbuf_size2_12_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_13_sram;
wire [0:1] mux_tree_tapbuf_size2_13_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_14_sram;
wire [0:1] mux_tree_tapbuf_size2_14_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_15_sram;
wire [0:1] mux_tree_tapbuf_size2_15_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_16_sram;
wire [0:1] mux_tree_tapbuf_size2_16_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_17_sram;
wire [0:1] mux_tree_tapbuf_size2_17_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_18_sram;
wire [0:1] mux_tree_tapbuf_size2_18_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_19_sram;
wire [0:1] mux_tree_tapbuf_size2_19_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_1_sram;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_20_sram;
wire [0:1] mux_tree_tapbuf_size2_20_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_21_sram;
wire [0:1] mux_tree_tapbuf_size2_21_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_22_sram;
wire [0:1] mux_tree_tapbuf_size2_22_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_23_sram;
wire [0:1] mux_tree_tapbuf_size2_23_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_24_sram;
wire [0:1] mux_tree_tapbuf_size2_24_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_25_sram;
wire [0:1] mux_tree_tapbuf_size2_25_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_26_sram;
wire [0:1] mux_tree_tapbuf_size2_26_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_2_sram;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_3_sram;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_4_sram;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_5_sram;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_6_sram;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_7_sram;
wire [0:1] mux_tree_tapbuf_size2_7_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_8_sram;
wire [0:1] mux_tree_tapbuf_size2_8_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_9_sram;
wire [0:1] mux_tree_tapbuf_size2_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_9_ccff_tail;
wire [0:1] mux_tree_tapbuf_size3_0_sram;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_10_sram;
wire [0:1] mux_tree_tapbuf_size3_10_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_11_sram;
wire [0:1] mux_tree_tapbuf_size3_11_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_12_sram;
wire [0:1] mux_tree_tapbuf_size3_12_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_13_sram;
wire [0:1] mux_tree_tapbuf_size3_13_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_14_sram;
wire [0:1] mux_tree_tapbuf_size3_14_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_15_sram;
wire [0:1] mux_tree_tapbuf_size3_15_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_16_sram;
wire [0:1] mux_tree_tapbuf_size3_16_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_17_sram;
wire [0:1] mux_tree_tapbuf_size3_17_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_18_sram;
wire [0:1] mux_tree_tapbuf_size3_18_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_19_sram;
wire [0:1] mux_tree_tapbuf_size3_19_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_1_sram;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_20_sram;
wire [0:1] mux_tree_tapbuf_size3_20_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_21_sram;
wire [0:1] mux_tree_tapbuf_size3_21_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_22_sram;
wire [0:1] mux_tree_tapbuf_size3_22_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_23_sram;
wire [0:1] mux_tree_tapbuf_size3_23_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_24_sram;
wire [0:1] mux_tree_tapbuf_size3_24_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_25_sram;
wire [0:1] mux_tree_tapbuf_size3_25_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_26_sram;
wire [0:1] mux_tree_tapbuf_size3_26_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_27_sram;
wire [0:1] mux_tree_tapbuf_size3_27_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_28_sram;
wire [0:1] mux_tree_tapbuf_size3_28_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_29_sram;
wire [0:1] mux_tree_tapbuf_size3_29_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_2_sram;
wire [0:1] mux_tree_tapbuf_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_30_sram;
wire [0:1] mux_tree_tapbuf_size3_30_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_31_sram;
wire [0:1] mux_tree_tapbuf_size3_31_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_32_sram;
wire [0:1] mux_tree_tapbuf_size3_32_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_33_sram;
wire [0:1] mux_tree_tapbuf_size3_33_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_34_sram;
wire [0:1] mux_tree_tapbuf_size3_34_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_35_sram;
wire [0:1] mux_tree_tapbuf_size3_35_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_36_sram;
wire [0:1] mux_tree_tapbuf_size3_36_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_37_sram;
wire [0:1] mux_tree_tapbuf_size3_37_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_38_sram;
wire [0:1] mux_tree_tapbuf_size3_38_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_39_sram;
wire [0:1] mux_tree_tapbuf_size3_39_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_3_sram;
wire [0:1] mux_tree_tapbuf_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_40_sram;
wire [0:1] mux_tree_tapbuf_size3_40_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_41_sram;
wire [0:1] mux_tree_tapbuf_size3_41_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_42_sram;
wire [0:1] mux_tree_tapbuf_size3_42_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_43_sram;
wire [0:1] mux_tree_tapbuf_size3_43_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_44_sram;
wire [0:1] mux_tree_tapbuf_size3_44_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_45_sram;
wire [0:1] mux_tree_tapbuf_size3_45_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_46_sram;
wire [0:1] mux_tree_tapbuf_size3_46_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_47_sram;
wire [0:1] mux_tree_tapbuf_size3_47_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_48_sram;
wire [0:1] mux_tree_tapbuf_size3_48_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_49_sram;
wire [0:1] mux_tree_tapbuf_size3_49_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_4_sram;
wire [0:1] mux_tree_tapbuf_size3_4_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_50_sram;
wire [0:1] mux_tree_tapbuf_size3_50_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_51_sram;
wire [0:1] mux_tree_tapbuf_size3_51_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_52_sram;
wire [0:1] mux_tree_tapbuf_size3_52_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_53_sram;
wire [0:1] mux_tree_tapbuf_size3_53_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_54_sram;
wire [0:1] mux_tree_tapbuf_size3_54_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_5_sram;
wire [0:1] mux_tree_tapbuf_size3_5_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_6_sram;
wire [0:1] mux_tree_tapbuf_size3_6_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_7_sram;
wire [0:1] mux_tree_tapbuf_size3_7_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_8_sram;
wire [0:1] mux_tree_tapbuf_size3_8_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_9_sram;
wire [0:1] mux_tree_tapbuf_size3_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size4_0_sram;
wire [0:2] mux_tree_tapbuf_size4_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_10_sram;
wire [0:2] mux_tree_tapbuf_size4_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_11_sram;
wire [0:2] mux_tree_tapbuf_size4_11_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_12_sram;
wire [0:2] mux_tree_tapbuf_size4_12_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_13_sram;
wire [0:2] mux_tree_tapbuf_size4_13_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_14_sram;
wire [0:2] mux_tree_tapbuf_size4_14_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_15_sram;
wire [0:2] mux_tree_tapbuf_size4_15_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_16_sram;
wire [0:2] mux_tree_tapbuf_size4_16_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_17_sram;
wire [0:2] mux_tree_tapbuf_size4_17_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_18_sram;
wire [0:2] mux_tree_tapbuf_size4_18_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_19_sram;
wire [0:2] mux_tree_tapbuf_size4_19_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_1_sram;
wire [0:2] mux_tree_tapbuf_size4_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_20_sram;
wire [0:2] mux_tree_tapbuf_size4_20_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_21_sram;
wire [0:2] mux_tree_tapbuf_size4_21_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_22_sram;
wire [0:2] mux_tree_tapbuf_size4_22_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_23_sram;
wire [0:2] mux_tree_tapbuf_size4_23_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_24_sram;
wire [0:2] mux_tree_tapbuf_size4_24_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_25_sram;
wire [0:2] mux_tree_tapbuf_size4_25_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_26_sram;
wire [0:2] mux_tree_tapbuf_size4_26_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_2_sram;
wire [0:2] mux_tree_tapbuf_size4_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_3_sram;
wire [0:2] mux_tree_tapbuf_size4_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_4_sram;
wire [0:2] mux_tree_tapbuf_size4_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_5_sram;
wire [0:2] mux_tree_tapbuf_size4_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_6_sram;
wire [0:2] mux_tree_tapbuf_size4_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_7_sram;
wire [0:2] mux_tree_tapbuf_size4_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_8_sram;
wire [0:2] mux_tree_tapbuf_size4_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_9_sram;
wire [0:2] mux_tree_tapbuf_size4_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size4_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size5_0_sram;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail;
wire [0:2] mux_tree_tapbuf_size7_0_sram;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_1_sram;
wire [0:2] mux_tree_tapbuf_size7_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_2_sram;
wire [0:2] mux_tree_tapbuf_size7_2_sram_inv;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_1_ccff_tail;
wire [0:3] mux_tree_tapbuf_size8_0_sram;
wire [0:3] mux_tree_tapbuf_size8_0_sram_inv;
wire [0:0] mux_tree_tapbuf_size8_mem_0_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[5] = chanx_right_in[4];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[7] = chanx_right_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[9] = chanx_right_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[57] = chanx_right_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[11] = chanx_right_in[10];
// ----- Local connection due to Wire 11 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[56] = chanx_right_in[11];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[13] = chanx_right_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[55] = chanx_right_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[15] = chanx_right_in[14];
// ----- Local connection due to Wire 15 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[54] = chanx_right_in[15];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[17] = chanx_right_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[53] = chanx_right_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[19] = chanx_right_in[18];
// ----- Local connection due to Wire 19 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[52] = chanx_right_in[19];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[23] = chanx_right_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[27] = chanx_right_in[26];
// ----- Local connection due to Wire 27 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[48] = chanx_right_in[27];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[47] = chanx_right_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[31] = chanx_right_in[30];
// ----- Local connection due to Wire 31 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[46] = chanx_right_in[31];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[33] = chanx_right_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[45] = chanx_right_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[35] = chanx_right_in[34];
// ----- Local connection due to Wire 35 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[44] = chanx_right_in[35];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[37] = chanx_right_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[43] = chanx_right_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[39] = chanx_right_in[38];
// ----- Local connection due to Wire 39 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[42] = chanx_right_in[39];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[41] = chanx_right_in[40];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[43] = chanx_right_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[45] = chanx_right_in[44];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[47] = chanx_right_in[46];
// ----- Local connection due to Wire 47 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[38] = chanx_right_in[47];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[49] = chanx_right_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[37] = chanx_right_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[51] = chanx_right_in[50];
// ----- Local connection due to Wire 51 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[36] = chanx_right_in[51];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[53] = chanx_right_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[35] = chanx_right_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[55] = chanx_right_in[54];
// ----- Local connection due to Wire 55 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[34] = chanx_right_in[55];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[57] = chanx_right_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[33] = chanx_right_in[57];
// ----- Local connection due to Wire 59 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[60] = chanx_right_in[59];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[61] = chanx_right_in[60];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[63] = chanx_right_in[62];
// ----- Local connection due to Wire 63 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[64] = chanx_right_in[63];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[5] = chanx_left_in[4];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[7] = chanx_left_in[6];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[9] = chanx_left_in[8];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[11] = chanx_left_in[10];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[13] = chanx_left_in[12];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[15] = chanx_left_in[14];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[17] = chanx_left_in[16];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[19] = chanx_left_in[18];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[23] = chanx_left_in[22];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[27] = chanx_left_in[26];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[31] = chanx_left_in[30];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[33] = chanx_left_in[32];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[35] = chanx_left_in[34];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[37] = chanx_left_in[36];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[39] = chanx_left_in[38];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[41] = chanx_left_in[40];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[43] = chanx_left_in[42];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[45] = chanx_left_in[44];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[47] = chanx_left_in[46];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[49] = chanx_left_in[48];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[51] = chanx_left_in[50];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[53] = chanx_left_in[52];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[55] = chanx_left_in[54];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[57] = chanx_left_in[56];
// ----- Local connection due to Wire 199 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[60] = chanx_left_in[59];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[61] = chanx_left_in[60];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[63] = chanx_left_in[62];
// ----- Local connection due to Wire 203 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[64] = chanx_left_in[63];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size3 mux_right_track_0 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[32]}),
		.sram(mux_tree_tapbuf_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_0_sram_inv[0:1]),
		.out(chanx_right_out[0]));

	mux_tree_tapbuf_size3 mux_right_track_2 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_, chany_bottom_in[31]}),
		.sram(mux_tree_tapbuf_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_1_sram_inv[0:1]),
		.out(chanx_right_out[1]));

	mux_tree_tapbuf_size3 mux_right_track_4 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[30], chany_bottom_in[64]}),
		.sram(mux_tree_tapbuf_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_2_sram_inv[0:1]),
		.out(chanx_right_out[2]));

	mux_tree_tapbuf_size3 mux_right_track_6 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, chany_bottom_in[29], chany_bottom_in[63]}),
		.sram(mux_tree_tapbuf_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_3_sram_inv[0:1]),
		.out(chanx_right_out[3]));

	mux_tree_tapbuf_size3 mux_right_track_28 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_, chany_bottom_in[23], chany_bottom_in[57]}),
		.sram(mux_tree_tapbuf_size3_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_4_sram_inv[0:1]),
		.out(chanx_right_out[14]));

	mux_tree_tapbuf_size3 mux_right_track_44 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[19], chany_bottom_in[53]}),
		.sram(mux_tree_tapbuf_size3_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_5_sram_inv[0:1]),
		.out(chanx_right_out[22]));

	mux_tree_tapbuf_size3 mux_right_track_48 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, chany_bottom_in[18], chany_bottom_in[52]}),
		.sram(mux_tree_tapbuf_size3_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_6_sram_inv[0:1]),
		.out(chanx_right_out[24]));

	mux_tree_tapbuf_size3 mux_right_track_52 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[17], chany_bottom_in[51]}),
		.sram(mux_tree_tapbuf_size3_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_7_sram_inv[0:1]),
		.out(chanx_right_out[26]));

	mux_tree_tapbuf_size3 mux_right_track_56 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, chany_bottom_in[16], chany_bottom_in[50]}),
		.sram(mux_tree_tapbuf_size3_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_8_sram_inv[0:1]),
		.out(chanx_right_out[28]));

	mux_tree_tapbuf_size3 mux_right_track_60 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[15], chany_bottom_in[49]}),
		.sram(mux_tree_tapbuf_size3_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_9_sram_inv[0:1]),
		.out(chanx_right_out[30]));

	mux_tree_tapbuf_size3 mux_right_track_64 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_, chany_bottom_in[14], chany_bottom_in[48]}),
		.sram(mux_tree_tapbuf_size3_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_10_sram_inv[0:1]),
		.out(chanx_right_out[32]));

	mux_tree_tapbuf_size3 mux_right_track_80 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[10], chany_bottom_in[44]}),
		.sram(mux_tree_tapbuf_size3_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_11_sram_inv[0:1]),
		.out(chanx_right_out[40]));

	mux_tree_tapbuf_size3 mux_right_track_84 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, chany_bottom_in[9], chany_bottom_in[43]}),
		.sram(mux_tree_tapbuf_size3_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_12_sram_inv[0:1]),
		.out(chanx_right_out[42]));

	mux_tree_tapbuf_size3 mux_right_track_88 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[8], chany_bottom_in[42]}),
		.sram(mux_tree_tapbuf_size3_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_13_sram_inv[0:1]),
		.out(chanx_right_out[44]));

	mux_tree_tapbuf_size3 mux_right_track_92 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, chany_bottom_in[7], chany_bottom_in[41]}),
		.sram(mux_tree_tapbuf_size3_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_14_sram_inv[0:1]),
		.out(chanx_right_out[46]));

	mux_tree_tapbuf_size3 mux_right_track_96 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[6], chany_bottom_in[40]}),
		.sram(mux_tree_tapbuf_size3_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_15_sram_inv[0:1]),
		.out(chanx_right_out[48]));

	mux_tree_tapbuf_size3 mux_right_track_100 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_, chany_bottom_in[5], chany_bottom_in[39]}),
		.sram(mux_tree_tapbuf_size3_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_16_sram_inv[0:1]),
		.out(chanx_right_out[50]));

	mux_tree_tapbuf_size3 mux_right_track_116 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[1], chany_bottom_in[35]}),
		.sram(mux_tree_tapbuf_size3_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_17_sram_inv[0:1]),
		.out(chanx_right_out[58]));

	mux_tree_tapbuf_size3 mux_bottom_track_17 (
		.in({chanx_right_in[20], chanx_left_in[15], chanx_left_in[20]}),
		.sram(mux_tree_tapbuf_size3_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_18_sram_inv[0:1]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_size3 mux_bottom_track_19 (
		.in({chanx_right_in[22], chanx_left_in[17], chanx_left_in[22]}),
		.sram(mux_tree_tapbuf_size3_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_19_sram_inv[0:1]),
		.out(chany_bottom_out[9]));

	mux_tree_tapbuf_size3 mux_bottom_track_21 (
		.in({chanx_right_in[24], chanx_left_in[19], chanx_left_in[24]}),
		.sram(mux_tree_tapbuf_size3_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_20_sram_inv[0:1]),
		.out(chany_bottom_out[10]));

	mux_tree_tapbuf_size3 mux_bottom_track_23 (
		.in({chanx_right_in[26], chanx_left_in[21], chanx_left_in[26]}),
		.sram(mux_tree_tapbuf_size3_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_21_sram_inv[0:1]),
		.out(chany_bottom_out[11]));

	mux_tree_tapbuf_size3 mux_bottom_track_25 (
		.in({chanx_right_in[28], chanx_left_in[23], chanx_left_in[28]}),
		.sram(mux_tree_tapbuf_size3_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_22_sram_inv[0:1]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_size3 mux_bottom_track_31 (
		.in({chanx_right_in[34], chanx_left_in[29], chanx_left_in[34]}),
		.sram(mux_tree_tapbuf_size3_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_23_sram_inv[0:1]),
		.out(chany_bottom_out[15]));

	mux_tree_tapbuf_size3 mux_bottom_track_33 (
		.in({chanx_right_in[36], chanx_left_in[31], chanx_left_in[36]}),
		.sram(mux_tree_tapbuf_size3_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_24_sram_inv[0:1]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_size3 mux_bottom_track_39 (
		.in({chanx_right_in[42], chanx_left_in[37], chanx_left_in[42]}),
		.sram(mux_tree_tapbuf_size3_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_25_sram_inv[0:1]),
		.out(chany_bottom_out[19]));

	mux_tree_tapbuf_size3 mux_bottom_track_41 (
		.in({chanx_right_in[44], chanx_left_in[39], chanx_left_in[44]}),
		.sram(mux_tree_tapbuf_size3_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_26_sram_inv[0:1]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_size3 mux_bottom_track_43 (
		.in({chanx_right_in[46], chanx_left_in[41], chanx_left_in[46]}),
		.sram(mux_tree_tapbuf_size3_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_27_sram_inv[0:1]),
		.out(chany_bottom_out[21]));

	mux_tree_tapbuf_size3 mux_bottom_track_49 (
		.in({chanx_right_in[52], chanx_left_in[47], chanx_left_in[52]}),
		.sram(mux_tree_tapbuf_size3_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_28_sram_inv[0:1]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_size3 mux_bottom_track_51 (
		.in({chanx_right_in[54], chanx_left_in[49], chanx_left_in[54]}),
		.sram(mux_tree_tapbuf_size3_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_29_sram_inv[0:1]),
		.out(chany_bottom_out[25]));

	mux_tree_tapbuf_size3 mux_bottom_track_53 (
		.in({chanx_right_in[56], chanx_left_in[51], chanx_left_in[56]}),
		.sram(mux_tree_tapbuf_size3_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_30_sram_inv[0:1]),
		.out(chany_bottom_out[26]));

	mux_tree_tapbuf_size3 mux_bottom_track_55 (
		.in({chanx_right_in[59], chanx_left_in[53], chanx_left_in[59]}),
		.sram(mux_tree_tapbuf_size3_31_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_31_sram_inv[0:1]),
		.out(chany_bottom_out[27]));

	mux_tree_tapbuf_size3 mux_bottom_track_63 (
		.in({chanx_right_in[61], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, chanx_left_in[61]}),
		.sram(mux_tree_tapbuf_size3_32_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_32_sram_inv[0:1]),
		.out(chany_bottom_out[31]));

	mux_tree_tapbuf_size3 mux_bottom_track_65 (
		.in({chanx_right_in[58], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, chanx_left_in[64]}),
		.sram(mux_tree_tapbuf_size3_33_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_33_sram_inv[0:1]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_size3 mux_bottom_track_81 (
		.in({chanx_right_in[43], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_}),
		.sram(mux_tree_tapbuf_size3_34_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_34_sram_inv[0:1]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_size3 mux_bottom_track_101 (
		.in({chanx_right_in[23], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_tree_tapbuf_size3_35_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_35_sram_inv[0:1]),
		.out(chany_bottom_out[50]));

	mux_tree_tapbuf_size3 mux_bottom_track_119 (
		.in({chanx_right_in[5], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_}),
		.sram(mux_tree_tapbuf_size3_36_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_36_sram_inv[0:1]),
		.out(chany_bottom_out[59]));

	mux_tree_tapbuf_size3 mux_bottom_track_125 (
		.in({chanx_right_in[1], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_}),
		.sram(mux_tree_tapbuf_size3_37_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_37_sram_inv[0:1]),
		.out(chany_bottom_out[62]));

	mux_tree_tapbuf_size3 mux_left_track_1 (
		.in({chany_bottom_in[33], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
		.sram(mux_tree_tapbuf_size3_38_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_38_sram_inv[0:1]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_size3 mux_left_track_5 (
		.in({chany_bottom_in[1], chany_bottom_in[35], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_39_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_39_sram_inv[0:1]),
		.out(chanx_left_out[2]));

	mux_tree_tapbuf_size3 mux_left_track_7 (
		.in({chany_bottom_in[2], chany_bottom_in[36], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_}),
		.sram(mux_tree_tapbuf_size3_40_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_40_sram_inv[0:1]),
		.out(chanx_left_out[3]));

	mux_tree_tapbuf_size3 mux_left_track_29 (
		.in({chany_bottom_in[8], chany_bottom_in[42], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
		.sram(mux_tree_tapbuf_size3_41_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_41_sram_inv[0:1]),
		.out(chanx_left_out[14]));

	mux_tree_tapbuf_size3 mux_left_track_45 (
		.in({chany_bottom_in[12], chany_bottom_in[46], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_42_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_42_sram_inv[0:1]),
		.out(chanx_left_out[22]));

	mux_tree_tapbuf_size3 mux_left_track_49 (
		.in({chany_bottom_in[13], chany_bottom_in[47], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size3_43_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_43_sram_inv[0:1]),
		.out(chanx_left_out[24]));

	mux_tree_tapbuf_size3 mux_left_track_53 (
		.in({chany_bottom_in[14], chany_bottom_in[48], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_44_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_44_sram_inv[0:1]),
		.out(chanx_left_out[26]));

	mux_tree_tapbuf_size3 mux_left_track_57 (
		.in({chany_bottom_in[15], chany_bottom_in[49], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_}),
		.sram(mux_tree_tapbuf_size3_45_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_45_sram_inv[0:1]),
		.out(chanx_left_out[28]));

	mux_tree_tapbuf_size3 mux_left_track_61 (
		.in({chany_bottom_in[16], chany_bottom_in[50], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
		.sram(mux_tree_tapbuf_size3_46_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_46_sram_inv[0:1]),
		.out(chanx_left_out[30]));

	mux_tree_tapbuf_size3 mux_left_track_65 (
		.in({chany_bottom_in[17], chany_bottom_in[51], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
		.sram(mux_tree_tapbuf_size3_47_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_47_sram_inv[0:1]),
		.out(chanx_left_out[32]));

	mux_tree_tapbuf_size3 mux_left_track_81 (
		.in({chany_bottom_in[21], chany_bottom_in[55], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_48_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_48_sram_inv[0:1]),
		.out(chanx_left_out[40]));

	mux_tree_tapbuf_size3 mux_left_track_85 (
		.in({chany_bottom_in[22], chany_bottom_in[56], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size3_49_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_49_sram_inv[0:1]),
		.out(chanx_left_out[42]));

	mux_tree_tapbuf_size3 mux_left_track_89 (
		.in({chany_bottom_in[23], chany_bottom_in[57], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_50_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_50_sram_inv[0:1]),
		.out(chanx_left_out[44]));

	mux_tree_tapbuf_size3 mux_left_track_93 (
		.in({chany_bottom_in[24], chany_bottom_in[58], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_}),
		.sram(mux_tree_tapbuf_size3_51_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_51_sram_inv[0:1]),
		.out(chanx_left_out[46]));

	mux_tree_tapbuf_size3 mux_left_track_97 (
		.in({chany_bottom_in[25], chany_bottom_in[59], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
		.sram(mux_tree_tapbuf_size3_52_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_52_sram_inv[0:1]),
		.out(chanx_left_out[48]));

	mux_tree_tapbuf_size3 mux_left_track_101 (
		.in({chany_bottom_in[26], chany_bottom_in[60], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
		.sram(mux_tree_tapbuf_size3_53_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_53_sram_inv[0:1]),
		.out(chanx_left_out[50]));

	mux_tree_tapbuf_size3 mux_left_track_117 (
		.in({chany_bottom_in[30], chany_bottom_in[64], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_54_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_54_sram_inv[0:1]),
		.out(chanx_left_out[58]));

	mux_tree_tapbuf_size3_mem mem_right_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size3_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_4_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_44 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_5_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_6_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_52 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_7_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_8_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_60 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_9_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_10_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_11_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_84 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_12_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_13_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_92 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_14_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_15_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_100 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_16_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_116 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_17_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_18_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_19_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_20_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_21_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_22_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_23_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_24_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_39 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_25_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_26_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_43 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_27_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_28_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_51 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_29_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_53 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_30_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_55 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_31_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_31_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_63 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_32_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_32_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_33_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_33_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_34_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_34_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_101 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_35_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_35_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_119 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_36_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_36_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_125 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_37_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_37_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_38_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_38_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_39_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_39_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_40_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_40_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_41_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_41_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_45 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_42_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_42_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_43_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_43_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_53 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_44_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_44_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_45_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_45_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_61 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_46_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_46_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_47_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_47_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_48_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_48_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_85 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_49_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_49_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_50_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_50_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_93 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_51_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_51_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_52_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_52_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_101 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_53_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_53_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_117 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_54_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_54_sram_inv[0:1]));

	mux_tree_tapbuf_size4 mux_right_track_8 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, chany_bottom_in[28], chany_bottom_in[62]}),
		.sram(mux_tree_tapbuf_size4_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_0_sram_inv[0:2]),
		.out(chanx_right_out[4]));

	mux_tree_tapbuf_size4 mux_right_track_12 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[27], chany_bottom_in[61]}),
		.sram(mux_tree_tapbuf_size4_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_1_sram_inv[0:2]),
		.out(chanx_right_out[6]));

	mux_tree_tapbuf_size4 mux_right_track_16 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, chany_bottom_in[26], chany_bottom_in[60]}),
		.sram(mux_tree_tapbuf_size4_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_2_sram_inv[0:2]),
		.out(chanx_right_out[8]));

	mux_tree_tapbuf_size4 mux_right_track_20 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[25], chany_bottom_in[59]}),
		.sram(mux_tree_tapbuf_size4_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_3_sram_inv[0:2]),
		.out(chanx_right_out[10]));

	mux_tree_tapbuf_size4 mux_right_track_24 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_, chany_bottom_in[24], chany_bottom_in[58]}),
		.sram(mux_tree_tapbuf_size4_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_4_sram_inv[0:2]),
		.out(chanx_right_out[12]));

	mux_tree_tapbuf_size4 mux_bottom_track_1 (
		.in({chanx_right_in[4], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, chanx_left_in[1], chanx_left_in[4]}),
		.sram(mux_tree_tapbuf_size4_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_5_sram_inv[0:2]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_size4 mux_bottom_track_3 (
		.in({chanx_right_in[6], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, chanx_left_in[2], chanx_left_in[6]}),
		.sram(mux_tree_tapbuf_size4_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_6_sram_inv[0:2]),
		.out(chany_bottom_out[1]));

	mux_tree_tapbuf_size4 mux_bottom_track_5 (
		.in({chanx_right_in[8], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[3], chanx_left_in[8]}),
		.sram(mux_tree_tapbuf_size4_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_7_sram_inv[0:2]),
		.out(chany_bottom_out[2]));

	mux_tree_tapbuf_size4 mux_bottom_track_7 (
		.in({chanx_right_in[10], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[5], chanx_left_in[10]}),
		.sram(mux_tree_tapbuf_size4_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_8_sram_inv[0:2]),
		.out(chany_bottom_out[3]));

	mux_tree_tapbuf_size4 mux_bottom_track_11 (
		.in({chanx_right_in[14], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, chanx_left_in[9], chanx_left_in[14]}),
		.sram(mux_tree_tapbuf_size4_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_9_sram_inv[0:2]),
		.out(chany_bottom_out[5]));

	mux_tree_tapbuf_size4 mux_bottom_track_13 (
		.in({chanx_right_in[16], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[11], chanx_left_in[16]}),
		.sram(mux_tree_tapbuf_size4_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_10_sram_inv[0:2]),
		.out(chany_bottom_out[6]));

	mux_tree_tapbuf_size4 mux_bottom_track_15 (
		.in({chanx_right_in[18], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[13], chanx_left_in[18]}),
		.sram(mux_tree_tapbuf_size4_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_11_sram_inv[0:2]),
		.out(chany_bottom_out[7]));

	mux_tree_tapbuf_size4 mux_bottom_track_27 (
		.in({chanx_right_in[30], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, chanx_left_in[25], chanx_left_in[30]}),
		.sram(mux_tree_tapbuf_size4_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_12_sram_inv[0:2]),
		.out(chany_bottom_out[13]));

	mux_tree_tapbuf_size4 mux_bottom_track_29 (
		.in({chanx_right_in[32], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, chanx_left_in[27], chanx_left_in[32]}),
		.sram(mux_tree_tapbuf_size4_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_13_sram_inv[0:2]),
		.out(chany_bottom_out[14]));

	mux_tree_tapbuf_size4 mux_bottom_track_35 (
		.in({chanx_right_in[38], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[33], chanx_left_in[38]}),
		.sram(mux_tree_tapbuf_size4_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_14_sram_inv[0:2]),
		.out(chany_bottom_out[17]));

	mux_tree_tapbuf_size4 mux_bottom_track_37 (
		.in({chanx_right_in[40], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[35], chanx_left_in[40]}),
		.sram(mux_tree_tapbuf_size4_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_15_sram_inv[0:2]),
		.out(chany_bottom_out[18]));

	mux_tree_tapbuf_size4 mux_bottom_track_45 (
		.in({chanx_right_in[48], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, chanx_left_in[43], chanx_left_in[48]}),
		.sram(mux_tree_tapbuf_size4_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_16_sram_inv[0:2]),
		.out(chany_bottom_out[22]));

	mux_tree_tapbuf_size4 mux_bottom_track_47 (
		.in({chanx_right_in[50], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, chanx_left_in[45], chanx_left_in[50]}),
		.sram(mux_tree_tapbuf_size4_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_17_sram_inv[0:2]),
		.out(chany_bottom_out[23]));

	mux_tree_tapbuf_size4 mux_bottom_track_57 (
		.in({chanx_right_in[60], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[55], chanx_left_in[60]}),
		.sram(mux_tree_tapbuf_size4_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_18_sram_inv[0:2]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_size4 mux_bottom_track_59 (
		.in({chanx_right_in[62], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[57], chanx_left_in[62]}),
		.sram(mux_tree_tapbuf_size4_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_19_sram_inv[0:2]),
		.out(chany_bottom_out[29]));

	mux_tree_tapbuf_size4 mux_bottom_track_61 (
		.in({chanx_right_in[63:64], chanx_left_in[58], chanx_left_in[63]}),
		.sram(mux_tree_tapbuf_size4_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_20_sram_inv[0:2]),
		.out(chany_bottom_out[30]));

	mux_tree_tapbuf_size4 mux_left_track_3 (
		.in({chany_bottom_in[0], chany_bottom_in[34], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
		.sram(mux_tree_tapbuf_size4_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_21_sram_inv[0:2]),
		.out(chanx_left_out[1]));

	mux_tree_tapbuf_size4 mux_left_track_9 (
		.in({chany_bottom_in[3], chany_bottom_in[37], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_size4_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_22_sram_inv[0:2]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_size4 mux_left_track_13 (
		.in({chany_bottom_in[4], chany_bottom_in[38], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size4_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_23_sram_inv[0:2]),
		.out(chanx_left_out[6]));

	mux_tree_tapbuf_size4 mux_left_track_17 (
		.in({chany_bottom_in[5], chany_bottom_in[39], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_}),
		.sram(mux_tree_tapbuf_size4_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_24_sram_inv[0:2]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_size4 mux_left_track_21 (
		.in({chany_bottom_in[6], chany_bottom_in[40], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
		.sram(mux_tree_tapbuf_size4_25_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_25_sram_inv[0:2]),
		.out(chanx_left_out[10]));

	mux_tree_tapbuf_size4 mux_left_track_25 (
		.in({chany_bottom_in[7], chany_bottom_in[41], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
		.sram(mux_tree_tapbuf_size4_26_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_26_sram_inv[0:2]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_size4_mem mem_right_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_0_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_right_track_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_1_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_right_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_2_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_right_track_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_3_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_right_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_4_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_5_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_6_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_7_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_8_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_9_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_10_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_11_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_12_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_13_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_35 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_14_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_37 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_15_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_45 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_16_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_47 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_17_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_18_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_59 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_19_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_61 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_20_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_21_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_22_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_23_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_24_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_25_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_25_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_26_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_26_sram_inv[0:2]));

	mux_tree_tapbuf_size2 mux_right_track_32 (
		.in({chany_bottom_in[22], chany_bottom_in[56]}),
		.sram(mux_tree_tapbuf_size2_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_0_sram_inv[0:1]),
		.out(chanx_right_out[16]));

	mux_tree_tapbuf_size2 mux_right_track_36 (
		.in({chany_bottom_in[21], chany_bottom_in[55]}),
		.sram(mux_tree_tapbuf_size2_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_1_sram_inv[0:1]),
		.out(chanx_right_out[18]));

	mux_tree_tapbuf_size2 mux_right_track_40 (
		.in({chany_bottom_in[20], chany_bottom_in[54]}),
		.sram(mux_tree_tapbuf_size2_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_2_sram_inv[0:1]),
		.out(chanx_right_out[20]));

	mux_tree_tapbuf_size2 mux_right_track_68 (
		.in({chany_bottom_in[13], chany_bottom_in[47]}),
		.sram(mux_tree_tapbuf_size2_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_3_sram_inv[0:1]),
		.out(chanx_right_out[34]));

	mux_tree_tapbuf_size2 mux_right_track_72 (
		.in({chany_bottom_in[12], chany_bottom_in[46]}),
		.sram(mux_tree_tapbuf_size2_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_4_sram_inv[0:1]),
		.out(chanx_right_out[36]));

	mux_tree_tapbuf_size2 mux_right_track_76 (
		.in({chany_bottom_in[11], chany_bottom_in[45]}),
		.sram(mux_tree_tapbuf_size2_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_5_sram_inv[0:1]),
		.out(chanx_right_out[38]));

	mux_tree_tapbuf_size2 mux_right_track_104 (
		.in({chany_bottom_in[4], chany_bottom_in[38]}),
		.sram(mux_tree_tapbuf_size2_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_6_sram_inv[0:1]),
		.out(chanx_right_out[52]));

	mux_tree_tapbuf_size2 mux_right_track_108 (
		.in({chany_bottom_in[3], chany_bottom_in[37]}),
		.sram(mux_tree_tapbuf_size2_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_7_sram_inv[0:1]),
		.out(chanx_right_out[54]));

	mux_tree_tapbuf_size2 mux_right_track_112 (
		.in({chany_bottom_in[2], chany_bottom_in[36]}),
		.sram(mux_tree_tapbuf_size2_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_8_sram_inv[0:1]),
		.out(chanx_right_out[56]));

	mux_tree_tapbuf_size2 mux_bottom_track_79 (
		.in({chanx_right_in[45], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_tree_tapbuf_size2_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_9_sram_inv[0:1]),
		.out(chany_bottom_out[39]));

	mux_tree_tapbuf_size2 mux_bottom_track_83 (
		.in({chanx_right_in[41], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_}),
		.sram(mux_tree_tapbuf_size2_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_10_sram_inv[0:1]),
		.out(chany_bottom_out[41]));

	mux_tree_tapbuf_size2 mux_bottom_track_99 (
		.in({chanx_right_in[25], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_}),
		.sram(mux_tree_tapbuf_size2_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_11_sram_inv[0:1]),
		.out(chany_bottom_out[49]));

	mux_tree_tapbuf_size2 mux_bottom_track_103 (
		.in({chanx_right_in[21], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_}),
		.sram(mux_tree_tapbuf_size2_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_12_sram_inv[0:1]),
		.out(chany_bottom_out[51]));

	mux_tree_tapbuf_size2 mux_bottom_track_117 (
		.in({chanx_right_in[7], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_}),
		.sram(mux_tree_tapbuf_size2_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_13_sram_inv[0:1]),
		.out(chany_bottom_out[58]));

	mux_tree_tapbuf_size2 mux_bottom_track_121 (
		.in({chanx_right_in[3], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_}),
		.sram(mux_tree_tapbuf_size2_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_14_sram_inv[0:1]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_size2 mux_bottom_track_123 (
		.in({chanx_right_in[2], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_tree_tapbuf_size2_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_15_sram_inv[0:1]),
		.out(chany_bottom_out[61]));

	mux_tree_tapbuf_size2 mux_bottom_track_127 (
		.in({chanx_right_in[0], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_}),
		.sram(mux_tree_tapbuf_size2_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_16_sram_inv[0:1]),
		.out(chany_bottom_out[63]));

	mux_tree_tapbuf_size2 mux_bottom_track_129 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, chanx_left_in[0]}),
		.sram(mux_tree_tapbuf_size2_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_17_sram_inv[0:1]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_size2 mux_left_track_33 (
		.in({chany_bottom_in[9], chany_bottom_in[43]}),
		.sram(mux_tree_tapbuf_size2_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_18_sram_inv[0:1]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_size2 mux_left_track_37 (
		.in({chany_bottom_in[10], chany_bottom_in[44]}),
		.sram(mux_tree_tapbuf_size2_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_19_sram_inv[0:1]),
		.out(chanx_left_out[18]));

	mux_tree_tapbuf_size2 mux_left_track_41 (
		.in({chany_bottom_in[11], chany_bottom_in[45]}),
		.sram(mux_tree_tapbuf_size2_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_20_sram_inv[0:1]),
		.out(chanx_left_out[20]));

	mux_tree_tapbuf_size2 mux_left_track_69 (
		.in({chany_bottom_in[18], chany_bottom_in[52]}),
		.sram(mux_tree_tapbuf_size2_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_21_sram_inv[0:1]),
		.out(chanx_left_out[34]));

	mux_tree_tapbuf_size2 mux_left_track_73 (
		.in({chany_bottom_in[19], chany_bottom_in[53]}),
		.sram(mux_tree_tapbuf_size2_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_22_sram_inv[0:1]),
		.out(chanx_left_out[36]));

	mux_tree_tapbuf_size2 mux_left_track_77 (
		.in({chany_bottom_in[20], chany_bottom_in[54]}),
		.sram(mux_tree_tapbuf_size2_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_23_sram_inv[0:1]),
		.out(chanx_left_out[38]));

	mux_tree_tapbuf_size2 mux_left_track_105 (
		.in({chany_bottom_in[27], chany_bottom_in[61]}),
		.sram(mux_tree_tapbuf_size2_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_24_sram_inv[0:1]),
		.out(chanx_left_out[52]));

	mux_tree_tapbuf_size2 mux_left_track_109 (
		.in({chany_bottom_in[28], chany_bottom_in[62]}),
		.sram(mux_tree_tapbuf_size2_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_25_sram_inv[0:1]),
		.out(chanx_left_out[54]));

	mux_tree_tapbuf_size2 mux_left_track_113 (
		.in({chany_bottom_in[29], chany_bottom_in[63]}),
		.sram(mux_tree_tapbuf_size2_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_26_sram_inv[0:1]),
		.out(chanx_left_out[56]));

	mux_tree_tapbuf_size2_mem mem_right_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_0_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_36 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_1_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_2_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_68 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_3_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_4_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_76 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_5_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_6_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_108 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_7_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_8_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_79 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_9_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_83 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_10_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_99 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_11_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_103 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_12_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_117 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_13_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_14_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_123 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_15_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_127 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_16_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_bottom_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_17_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_18_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_37 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_19_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_20_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_69 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_21_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_22_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_77 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_23_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_24_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_109 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_25_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_26_sram_inv[0:1]));

	mux_tree_tapbuf_size8 mux_right_track_118 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_, chany_bottom_in[0], chany_bottom_in[34]}),
		.sram(mux_tree_tapbuf_size8_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_0_sram_inv[0:3]),
		.out(chanx_right_out[59]));

	mux_tree_tapbuf_size8_mem mem_right_track_118 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_0_sram_inv[0:3]));

	mux_tree_tapbuf_size7 mux_right_track_124 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_, chany_bottom_in[33]}),
		.sram(mux_tree_tapbuf_size7_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_0_sram_inv[0:2]),
		.out(chanx_right_out[62]));

	mux_tree_tapbuf_size7 mux_left_track_119 (
		.in({chany_bottom_in[31], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
		.sram(mux_tree_tapbuf_size7_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_1_sram_inv[0:2]),
		.out(chanx_left_out[59]));

	mux_tree_tapbuf_size7 mux_left_track_125 (
		.in({chany_bottom_in[32], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
		.sram(mux_tree_tapbuf_size7_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_2_sram_inv[0:2]),
		.out(chanx_left_out[62]));

	mux_tree_tapbuf_size7_mem mem_right_track_124 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_0_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_119 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_1_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_125 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_1_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_2_sram_inv[0:2]));

	mux_tree_tapbuf_size5 mux_bottom_track_9 (
		.in({chanx_right_in[12], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, chanx_left_in[7], chanx_left_in[12]}),
		.sram(mux_tree_tapbuf_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_0_sram_inv[0:2]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_0_sram_inv[0:2]));

endmodule
// ----- END Verilog module for sb_1__4_ -----

//----- Default net type -----
`default_nettype wire



