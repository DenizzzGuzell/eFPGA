//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Tile Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed Aug 14 09:11:37 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype wire

// ----- Verilog module for tile_1__5_ -----
module tile_1__5_(prog_clk,
                  sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
                  sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_,
                  sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                  sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_,
                  sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
                  sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_,
                  sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_,
                  sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_,
                  sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_,
                  sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_,
                  sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
                  sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_,
                  sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                  sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_,
                  sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
                  sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_,
                  sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
                  sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_,
                  sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                  sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_,
                  sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
                  sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_,
                  sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_,
                  sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_,
                  sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_,
                  sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_,
                  sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
                  sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_,
                  sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                  sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_,
                  sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
                  sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_,
                  sb_1__4__chany_bottom_in,
                  sb_2__4__chanx_right_in,
                  sb_2__4__chany_bottom_in,
                  grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_,
                  grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_,
                  grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_,
                  grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_,
                  grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_,
                  grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_,
                  grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_,
                  grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_,
                  grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_,
                  cbx_1__4__chanx_left_in,
                  cby_2__5__chany_top_in,
                  ccff_head,
                  cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_,
                  cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_,
                  cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_,
                  cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_,
                  cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_,
                  cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_,
                  cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_,
                  cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_,
                  cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_,
                  cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_,
                  cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_,
                  cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_,
                  cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_,
                  cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_,
                  cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_,
                  cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_,
                  cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_,
                  cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_,
                  cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_,
                  cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_,
                  cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_,
                  cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_,
                  cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_,
                  cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_,
                  sb_1__4__chany_bottom_out,
                  sb_2__4__chanx_right_out,
                  sb_2__4__chany_bottom_out,
                  grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_,
                  grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_,
                  grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_,
                  grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_,
                  grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_,
                  grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_,
                  grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_,
                  grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_,
                  cbx_1__4__chanx_left_out,
                  cby_2__5__chany_top_out,
                  ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
//----- INPUT PORTS -----
input [0:0] sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_;
//----- INPUT PORTS -----
input [0:0] sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
//----- INPUT PORTS -----
input [0:0] sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
//----- INPUT PORTS -----
input [0:0] sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
//----- INPUT PORTS -----
input [0:0] sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
//----- INPUT PORTS -----
input [0:0] sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
//----- INPUT PORTS -----
input [0:0] sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_;
//----- INPUT PORTS -----
input [0:0] sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
//----- INPUT PORTS -----
input [0:0] sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_;
//----- INPUT PORTS -----
input [0:0] sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
//----- INPUT PORTS -----
input [0:0] sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
//----- INPUT PORTS -----
input [0:0] sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
//----- INPUT PORTS -----
input [0:0] sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
//----- INPUT PORTS -----
input [0:0] sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
//----- INPUT PORTS -----
input [0:0] sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_;
//----- INPUT PORTS -----
input [0:64] sb_1__4__chany_bottom_in;
//----- INPUT PORTS -----
input [0:64] sb_2__4__chanx_right_in;
//----- INPUT PORTS -----
input [0:64] sb_2__4__chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_;
//----- INPUT PORTS -----
input [0:0] grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_;
//----- INPUT PORTS -----
input [0:0] grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_;
//----- INPUT PORTS -----
input [0:0] grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_;
//----- INPUT PORTS -----
input [0:0] grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_;
//----- INPUT PORTS -----
input [0:0] grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_;
//----- INPUT PORTS -----
input [0:0] grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_;
//----- INPUT PORTS -----
input [0:0] grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_;
//----- INPUT PORTS -----
input [0:0] grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_;
//----- INPUT PORTS -----
input [0:64] cbx_1__4__chanx_left_in;
//----- INPUT PORTS -----
input [0:64] cby_2__5__chany_top_in;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
//----- OUTPUT PORTS -----
output [0:64] sb_1__4__chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:64] sb_2__4__chanx_right_out;
//----- OUTPUT PORTS -----
output [0:64] sb_2__4__chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:0] grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
//----- OUTPUT PORTS -----
output [0:0] grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
//----- OUTPUT PORTS -----
output [0:0] grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
//----- OUTPUT PORTS -----
output [0:0] grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
//----- OUTPUT PORTS -----
output [0:0] grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
//----- OUTPUT PORTS -----
output [0:0] grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
//----- OUTPUT PORTS -----
output [0:0] grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
//----- OUTPUT PORTS -----
output [0:0] grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
//----- OUTPUT PORTS -----
output [0:64] cbx_1__4__chanx_left_out;
//----- OUTPUT PORTS -----
output [0:64] cby_2__5__chany_top_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:0] cbx_1__4__0_ccff_tail;
wire [0:64] cbx_1__4__0_chanx_right_out;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_0_;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_1_;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_2_;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_3_;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_4_;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_5_;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_6_;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_7_;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_8_;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_9_;
wire [0:0] cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cbx_1__9__0_ccff_tail;
wire [0:64] cbx_1__9__0_chanx_left_out;
wire [0:64] cbx_1__9__0_chanx_right_out;
wire [0:64] cby_2__5__0_chany_bottom_out;
wire [0:0] sb_1__4__0_ccff_tail;
wire [0:64] sb_1__4__0_chanx_left_out;
wire [0:64] sb_1__4__0_chanx_right_out;
wire [0:64] sb_2__4__0_chanx_left_out;
wire [0:64] sb_2__4__0_chany_top_out;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	grid_memory grid_memory_1__5_ (
		.top_width_0_height_0_subtile_0__pin_d_in_0_(grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.top_width_0_height_0_subtile_0__pin_d_in_1_(grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.top_width_0_height_0_subtile_0__pin_d_in_2_(grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.top_width_0_height_0_subtile_0__pin_d_in_3_(grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.top_width_0_height_0_subtile_0__pin_d_in_4_(grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.top_width_0_height_0_subtile_0__pin_d_in_5_(grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.top_width_0_height_0_subtile_0__pin_d_in_6_(grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.top_width_0_height_0_subtile_0__pin_d_in_7_(grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.bottom_width_0_height_0_subtile_0__pin_addr_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_0_),
		.bottom_width_0_height_0_subtile_0__pin_addr_1_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_1_),
		.bottom_width_0_height_0_subtile_0__pin_addr_2_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_2_),
		.bottom_width_0_height_0_subtile_0__pin_addr_3_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_3_),
		.bottom_width_0_height_0_subtile_0__pin_addr_4_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_4_),
		.bottom_width_0_height_0_subtile_0__pin_addr_5_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_5_),
		.bottom_width_0_height_0_subtile_0__pin_addr_6_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_6_),
		.bottom_width_0_height_0_subtile_0__pin_addr_7_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_7_),
		.bottom_width_0_height_0_subtile_0__pin_addr_8_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_8_),
		.bottom_width_0_height_0_subtile_0__pin_addr_9_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_9_),
		.bottom_width_0_height_0_subtile_0__pin_wen_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_wen_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_),
		.top_width_0_height_0_subtile_0__pin_d_out_0_(grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.top_width_0_height_0_subtile_0__pin_d_out_1_(grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.top_width_0_height_0_subtile_0__pin_d_out_2_(grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.top_width_0_height_0_subtile_0__pin_d_out_3_(grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.top_width_0_height_0_subtile_0__pin_d_out_4_(grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.top_width_0_height_0_subtile_0__pin_d_out_5_(grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.top_width_0_height_0_subtile_0__pin_d_out_6_(grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.top_width_0_height_0_subtile_0__pin_d_out_7_(grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_));

	cbx_1__4_ cbx_1__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_1__4__chanx_left_in[0:64]),
		.chanx_right_in(sb_1__4__0_chanx_left_out[0:64]),
		.ccff_head(ccff_head),
		.chanx_left_out(cbx_1__4__chanx_left_out[0:64]),
		.chanx_right_out(cbx_1__4__0_chanx_right_out[0:64]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_addr_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_addr_1_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_addr_2_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_addr_3_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_addr_4_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_addr_5_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_addr_6_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_addr_7_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_addr_8_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_addr_9_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_addr_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_wen_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.ccff_tail(cbx_1__4__0_ccff_tail));

	cbx_1__9_ cbx_2__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__0_chanx_right_out[0:64]),
		.chanx_right_in(sb_2__4__0_chanx_left_out[0:64]),
		.ccff_head(cbx_1__4__0_ccff_tail),
		.chanx_left_out(cbx_1__9__0_chanx_left_out[0:64]),
		.chanx_right_out(cbx_1__9__0_chanx_right_out[0:64]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_2__4__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.ccff_tail(cbx_1__9__0_ccff_tail));

	cby_2__5_ cby_2__5_ (
		.chany_bottom_in(sb_2__4__0_chany_top_out[0:64]),
		.chany_top_in(cby_2__5__chany_top_in[0:64]),
		.chany_bottom_out(cby_2__5__0_chany_bottom_out[0:64]),
		.chany_top_out(cby_2__5__chany_top_out[0:64]));

	sb_1__4_ sb_1__4_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__9__0_chanx_left_out[0:64]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(sb_1__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_),
		.chany_bottom_in(sb_1__4__chany_bottom_in[0:64]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_1__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__4__0_chanx_right_out[0:64]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(sb_1__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_),
		.ccff_head(cbx_1__9__0_ccff_tail),
		.chanx_right_out(sb_1__4__0_chanx_right_out[0:64]),
		.chany_bottom_out(sb_1__4__chany_bottom_out[0:64]),
		.chanx_left_out(sb_1__4__0_chanx_left_out[0:64]),
		.ccff_tail(sb_1__4__0_ccff_tail));

	sb_2__4_ sb_2__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_2__5__0_chany_bottom_out[0:64]),
		.chanx_right_in(sb_2__4__chanx_right_in[0:64]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(sb_2__4__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_),
		.chany_bottom_in(sb_2__4__chany_bottom_in[0:64]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_2__4__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__9__0_chanx_right_out[0:64]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(sb_2__4__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_),
		.ccff_head(sb_1__4__0_ccff_tail),
		.chany_top_out(sb_2__4__0_chany_top_out[0:64]),
		.chanx_right_out(sb_2__4__chanx_right_out[0:64]),
		.chany_bottom_out(sb_2__4__chany_bottom_out[0:64]),
		.chanx_left_out(sb_2__4__0_chanx_left_out[0:64]),
		.ccff_tail(ccff_tail));

endmodule
// ----- END Verilog module for tile_1__5_ -----

//----- Default net type -----
`default_nettype wire




