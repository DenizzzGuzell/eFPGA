//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Top-level Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Tue Jul 30 05:35:22 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype wire

// ----- Verilog module for fpga_top -----
module _fpga_top(clk,
                Reset,
                prog_clk,
                IO_ISOL_N,
                gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN,
                gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT,
                gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR,
                ccff_head,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] clk;
//----- GLOBAL PORTS -----
input [0:0] Reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- GLOBAL PORTS -----
input [0:0] IO_ISOL_N;
//----- GPIN PORTS -----
input [0:63] gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN;
//----- GPOUT PORTS -----
output [0:63] gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT;
//----- GPOUT PORTS -----
output [0:63] gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR;
//----- INPUT PORTS -----
input [0:31] ccff_head;
//----- OUTPUT PORTS -----
output [0:31] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:0] direct_interc_0_out;
wire [0:0] direct_interc_10_out;
wire [0:0] direct_interc_11_out;
wire [0:0] direct_interc_12_out;
wire [0:0] direct_interc_13_out;
wire [0:0] direct_interc_14_out;
wire [0:0] direct_interc_15_out;
wire [0:0] direct_interc_16_out;
wire [0:0] direct_interc_17_out;
wire [0:0] direct_interc_18_out;
wire [0:0] direct_interc_19_out;
wire [0:0] direct_interc_1_out;
wire [0:0] direct_interc_20_out;
wire [0:0] direct_interc_21_out;
wire [0:0] direct_interc_22_out;
wire [0:0] direct_interc_23_out;
wire [0:0] direct_interc_24_out;
wire [0:0] direct_interc_25_out;
wire [0:0] direct_interc_26_out;
wire [0:0] direct_interc_27_out;
wire [0:0] direct_interc_2_out;
wire [0:0] direct_interc_3_out;
wire [0:0] direct_interc_4_out;
wire [0:0] direct_interc_5_out;
wire [0:0] direct_interc_6_out;
wire [0:0] direct_interc_7_out;
wire [0:0] direct_interc_8_out;
wire [0:0] direct_interc_9_out;
wire [0:64] tile_0__1__0_cby_0__1__chany_top_out;
wire [0:0] tile_0__1__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__1__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__1__0_sb_0__0__chanx_right_out;
wire [0:64] tile_0__2__0_cby_0__2__chany_top_out;
wire [0:0] tile_0__2__0_ccff_tail;
wire [0:0] tile_0__2__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__2__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__2__0_sb_0__1__chanx_right_out;
wire [0:64] tile_0__2__0_sb_0__1__chany_bottom_out;
wire [0:64] tile_0__2__1_cby_0__2__chany_top_out;
wire [0:0] tile_0__2__1_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__2__1_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__2__1_sb_0__1__chanx_right_out;
wire [0:64] tile_0__2__1_sb_0__1__chany_bottom_out;
wire [0:64] tile_0__2__2_cby_0__2__chany_top_out;
wire [0:0] tile_0__2__2_ccff_tail;
wire [0:0] tile_0__2__2_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__2__2_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__2__2_sb_0__1__chanx_right_out;
wire [0:64] tile_0__2__2_sb_0__1__chany_bottom_out;
wire [0:64] tile_0__2__3_cby_0__2__chany_top_out;
wire [0:0] tile_0__2__3_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__2__3_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__2__3_sb_0__1__chanx_right_out;
wire [0:64] tile_0__2__3_sb_0__1__chany_bottom_out;
wire [0:64] tile_0__2__4_cby_0__2__chany_top_out;
wire [0:0] tile_0__2__4_ccff_tail;
wire [0:0] tile_0__2__4_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__2__4_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__2__4_sb_0__1__chanx_right_out;
wire [0:64] tile_0__2__4_sb_0__1__chany_bottom_out;
wire [0:64] tile_0__2__5_cby_0__2__chany_top_out;
wire [0:0] tile_0__2__5_ccff_tail;
wire [0:0] tile_0__2__5_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__2__5_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__2__5_sb_0__1__chanx_right_out;
wire [0:64] tile_0__2__5_sb_0__1__chany_bottom_out;
wire [0:64] tile_0__2__6_cby_0__2__chany_top_out;
wire [0:0] tile_0__2__6_ccff_tail;
wire [0:0] tile_0__2__6_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_0__2__6_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_0__2__6_sb_0__1__chanx_right_out;
wire [0:64] tile_0__2__6_sb_0__1__chany_bottom_out;
wire [0:64] tile_0__9__0_sb_0__8__chanx_right_out;
wire [0:64] tile_0__9__0_sb_0__8__chany_bottom_out;
wire [0:0] tile_1__0__0_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__0_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__1_ccff_tail;
wire [0:0] tile_1__0__1_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__1_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__2_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__2_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__3_ccff_tail;
wire [0:0] tile_1__0__3_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__3_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__4_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__4_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__5_ccff_tail;
wire [0:0] tile_1__0__5_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__5_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__6_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__6_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__0__7_ccff_tail;
wire [0:0] tile_1__0__7_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__0__7_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_1__1__0_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_1__1__0_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_1__1__0_cbx_1__0__chanx_left_out;
wire [0:64] tile_1__1__0_cby_1__1__chany_top_out;
wire [0:0] tile_1__1__0_ccff_tail;
wire [0:0] tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__1__0_sb_1__0__chanx_right_out;
wire [0:0] tile_1__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__0_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__0_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__0_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__0_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__1_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__1_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__1_ccff_tail;
wire [0:0] tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__1_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__1_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__2_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__2_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__2_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__2_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__3_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__3_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__3_ccff_tail;
wire [0:0] tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__3_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__3_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__4_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__4_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__4_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__4_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__5_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__5_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__5_ccff_tail;
wire [0:0] tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__5_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__5_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__2__6_cbx_1__1__chanx_left_out;
wire [0:64] tile_1__2__6_cby_1__2__chany_top_out;
wire [0:0] tile_1__2__6_ccff_tail;
wire [0:0] tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_1__2__6_sb_1__1__chanx_right_out;
wire [0:64] tile_1__2__6_sb_1__1__chany_bottom_out;
wire [0:0] tile_1__8__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_1__9__0_cbx_1__8__chanx_left_out;
wire [0:0] tile_1__9__0_ccff_tail;
wire [0:0] tile_1__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_1__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_1__9__0_sb_1__8__chanx_right_out;
wire [0:64] tile_1__9__0_sb_1__8__chany_bottom_out;
wire [0:0] tile_2__1__0_cbx_2__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_2__1__0_cbx_2__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_2__1__0_cbx_2__0__chanx_left_out;
wire [0:0] tile_2__1__0_cbx_3__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_2__1__0_cbx_3__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_2__1__0_cby_3__1__chany_top_out;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_;
wire [0:64] tile_2__1__0_sb_3__0__chanx_right_out;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_;
wire [0:0] tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_;
wire [0:64] tile_2__2__0_cbx_2__1__chanx_left_out;
wire [0:64] tile_2__2__0_cby_3__2__chany_top_out;
wire [0:0] tile_2__2__0_ccff_tail;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_;
wire [0:64] tile_2__2__0_sb_3__1__chanx_right_out;
wire [0:64] tile_2__2__0_sb_3__1__chany_bottom_out;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_;
wire [0:0] tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_;
wire [0:64] tile_2__2__1_cbx_2__1__chanx_left_out;
wire [0:64] tile_2__2__1_cby_3__2__chany_top_out;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_;
wire [0:64] tile_2__2__1_sb_3__1__chanx_right_out;
wire [0:64] tile_2__2__1_sb_3__1__chany_bottom_out;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_;
wire [0:0] tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_;
wire [0:64] tile_2__2__2_cbx_2__1__chanx_left_out;
wire [0:64] tile_2__2__2_cby_3__2__chany_top_out;
wire [0:0] tile_2__2__2_ccff_tail;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_;
wire [0:64] tile_2__2__2_sb_3__1__chanx_right_out;
wire [0:64] tile_2__2__2_sb_3__1__chany_bottom_out;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_;
wire [0:0] tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_;
wire [0:64] tile_2__2__3_cbx_2__1__chanx_left_out;
wire [0:64] tile_2__2__3_cby_3__2__chany_top_out;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_;
wire [0:64] tile_2__2__3_sb_3__1__chanx_right_out;
wire [0:64] tile_2__2__3_sb_3__1__chany_bottom_out;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_;
wire [0:0] tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_;
wire [0:64] tile_2__2__4_cbx_2__1__chanx_left_out;
wire [0:64] tile_2__2__4_cby_3__2__chany_top_out;
wire [0:0] tile_2__2__4_ccff_tail;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_;
wire [0:64] tile_2__2__4_sb_3__1__chanx_right_out;
wire [0:64] tile_2__2__4_sb_3__1__chany_bottom_out;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_;
wire [0:0] tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_;
wire [0:64] tile_2__2__5_cbx_2__1__chanx_left_out;
wire [0:64] tile_2__2__5_cby_3__2__chany_top_out;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_;
wire [0:64] tile_2__2__5_sb_3__1__chanx_right_out;
wire [0:64] tile_2__2__5_sb_3__1__chany_bottom_out;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_;
wire [0:0] tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_;
wire [0:64] tile_2__2__6_cbx_2__1__chanx_left_out;
wire [0:64] tile_2__2__6_cby_3__2__chany_top_out;
wire [0:0] tile_2__2__6_ccff_tail;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_;
wire [0:0] tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_;
wire [0:64] tile_2__2__6_sb_3__1__chanx_right_out;
wire [0:64] tile_2__2__6_sb_3__1__chany_bottom_out;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_;
wire [0:0] tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_;
wire [0:64] tile_2__9__0_cbx_2__8__chanx_left_out;
wire [0:0] tile_2__9__0_ccff_tail;
wire [0:0] tile_2__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_2__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_2__9__0_sb_2__8__chanx_right_out;
wire [0:64] tile_3__9__0_cbx_3__8__chanx_left_out;
wire [0:0] tile_3__9__0_ccff_tail;
wire [0:0] tile_3__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_3__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_3__9__0_sb_3__8__chanx_right_out;
wire [0:64] tile_3__9__0_sb_3__8__chany_bottom_out;
wire [0:0] tile_4__1__0_cbx_4__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_4__1__0_cbx_4__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_4__1__0_cbx_4__0__chanx_left_out;
wire [0:64] tile_4__1__0_cby_4__1__chany_top_out;
wire [0:0] tile_4__1__0_ccff_tail;
wire [0:0] tile_4__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_4__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_4__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_4__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_4__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_4__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_4__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_4__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_4__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_4__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_4__1__0_sb_4__0__chanx_right_out;
wire [0:0] tile_4__1__1_cbx_4__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_4__1__1_cbx_4__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_4__1__1_cbx_4__0__chanx_left_out;
wire [0:64] tile_4__1__1_cby_4__1__chany_top_out;
wire [0:0] tile_4__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_4__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_4__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_4__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_4__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_4__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_4__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_4__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_4__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_4__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_4__1__1_sb_4__0__chanx_right_out;
wire [0:0] tile_4__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_4__2__0_cbx_4__1__chanx_left_out;
wire [0:64] tile_4__2__0_cby_4__2__chany_top_out;
wire [0:0] tile_4__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_4__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_4__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_4__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_4__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_4__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_4__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_4__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_4__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_4__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_4__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_4__2__0_sb_4__1__chanx_right_out;
wire [0:64] tile_4__2__0_sb_4__1__chany_bottom_out;
wire [0:0] tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_4__2__10_cbx_4__1__chanx_left_out;
wire [0:64] tile_4__2__10_cby_4__2__chany_top_out;
wire [0:0] tile_4__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_4__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_4__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_4__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_4__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_4__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_4__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_4__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_4__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_4__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_4__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_4__2__10_sb_4__1__chanx_right_out;
wire [0:64] tile_4__2__10_sb_4__1__chany_bottom_out;
wire [0:0] tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_4__2__11_cbx_4__1__chanx_left_out;
wire [0:64] tile_4__2__11_cby_4__2__chany_top_out;
wire [0:0] tile_4__2__11_ccff_tail;
wire [0:0] tile_4__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_4__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_4__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_4__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_4__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_4__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_4__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_4__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_4__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_4__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_4__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_4__2__11_sb_4__1__chanx_right_out;
wire [0:64] tile_4__2__11_sb_4__1__chany_bottom_out;
wire [0:0] tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_4__2__12_cbx_4__1__chanx_left_out;
wire [0:64] tile_4__2__12_cby_4__2__chany_top_out;
wire [0:0] tile_4__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_4__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_4__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_4__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_4__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_4__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_4__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_4__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_4__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_4__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_4__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_4__2__12_sb_4__1__chanx_right_out;
wire [0:64] tile_4__2__12_sb_4__1__chany_bottom_out;
wire [0:0] tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_4__2__13_cbx_4__1__chanx_left_out;
wire [0:64] tile_4__2__13_cby_4__2__chany_top_out;
wire [0:0] tile_4__2__13_ccff_tail;
wire [0:0] tile_4__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_4__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_4__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_4__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_4__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_4__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_4__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_4__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_4__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_4__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_4__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_4__2__13_sb_4__1__chanx_right_out;
wire [0:64] tile_4__2__13_sb_4__1__chany_bottom_out;
wire [0:0] tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_4__2__1_cbx_4__1__chanx_left_out;
wire [0:64] tile_4__2__1_cby_4__2__chany_top_out;
wire [0:0] tile_4__2__1_ccff_tail;
wire [0:0] tile_4__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_4__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_4__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_4__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_4__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_4__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_4__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_4__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_4__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_4__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_4__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_4__2__1_sb_4__1__chanx_right_out;
wire [0:64] tile_4__2__1_sb_4__1__chany_bottom_out;
wire [0:0] tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_4__2__2_cbx_4__1__chanx_left_out;
wire [0:64] tile_4__2__2_cby_4__2__chany_top_out;
wire [0:0] tile_4__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_4__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_4__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_4__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_4__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_4__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_4__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_4__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_4__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_4__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_4__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_4__2__2_sb_4__1__chanx_right_out;
wire [0:64] tile_4__2__2_sb_4__1__chany_bottom_out;
wire [0:0] tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_4__2__3_cbx_4__1__chanx_left_out;
wire [0:64] tile_4__2__3_cby_4__2__chany_top_out;
wire [0:0] tile_4__2__3_ccff_tail;
wire [0:0] tile_4__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_4__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_4__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_4__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_4__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_4__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_4__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_4__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_4__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_4__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_4__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_4__2__3_sb_4__1__chanx_right_out;
wire [0:64] tile_4__2__3_sb_4__1__chany_bottom_out;
wire [0:0] tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_4__2__4_cbx_4__1__chanx_left_out;
wire [0:64] tile_4__2__4_cby_4__2__chany_top_out;
wire [0:0] tile_4__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_4__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_4__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_4__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_4__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_4__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_4__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_4__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_4__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_4__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_4__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_4__2__4_sb_4__1__chanx_right_out;
wire [0:64] tile_4__2__4_sb_4__1__chany_bottom_out;
wire [0:0] tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_4__2__5_cbx_4__1__chanx_left_out;
wire [0:64] tile_4__2__5_cby_4__2__chany_top_out;
wire [0:0] tile_4__2__5_ccff_tail;
wire [0:0] tile_4__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_4__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_4__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_4__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_4__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_4__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_4__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_4__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_4__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_4__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_4__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_4__2__5_sb_4__1__chanx_right_out;
wire [0:64] tile_4__2__5_sb_4__1__chany_bottom_out;
wire [0:0] tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_4__2__6_cbx_4__1__chanx_left_out;
wire [0:64] tile_4__2__6_cby_4__2__chany_top_out;
wire [0:0] tile_4__2__6_ccff_tail;
wire [0:0] tile_4__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_4__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_4__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_4__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_4__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_4__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_4__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_4__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_4__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_4__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_4__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_4__2__6_sb_4__1__chanx_right_out;
wire [0:64] tile_4__2__6_sb_4__1__chany_bottom_out;
wire [0:0] tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_4__2__7_cbx_4__1__chanx_left_out;
wire [0:64] tile_4__2__7_cby_4__2__chany_top_out;
wire [0:0] tile_4__2__7_ccff_tail;
wire [0:0] tile_4__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_4__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_4__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_4__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_4__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_4__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_4__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_4__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_4__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_4__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_4__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_4__2__7_sb_4__1__chanx_right_out;
wire [0:64] tile_4__2__7_sb_4__1__chany_bottom_out;
wire [0:0] tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_4__2__8_cbx_4__1__chanx_left_out;
wire [0:64] tile_4__2__8_cby_4__2__chany_top_out;
wire [0:0] tile_4__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_4__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_4__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_4__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_4__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_4__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_4__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_4__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_4__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_4__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_4__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_4__2__8_sb_4__1__chanx_right_out;
wire [0:64] tile_4__2__8_sb_4__1__chany_bottom_out;
wire [0:0] tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_4__2__9_cbx_4__1__chanx_left_out;
wire [0:64] tile_4__2__9_cby_4__2__chany_top_out;
wire [0:0] tile_4__2__9_ccff_tail;
wire [0:0] tile_4__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_4__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_4__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_4__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_4__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_4__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_4__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_4__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_4__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_4__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_4__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_4__2__9_sb_4__1__chanx_right_out;
wire [0:64] tile_4__2__9_sb_4__1__chany_bottom_out;
wire [0:0] tile_4__8__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_4__9__0_cbx_4__8__chanx_left_out;
wire [0:0] tile_4__9__0_ccff_tail;
wire [0:0] tile_4__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_4__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_4__9__0_sb_4__8__chanx_right_out;
wire [0:64] tile_4__9__0_sb_4__8__chany_bottom_out;
wire [0:0] tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_4__9__1_cbx_4__8__chanx_left_out;
wire [0:0] tile_4__9__1_ccff_tail;
wire [0:0] tile_4__9__1_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_4__9__1_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_4__9__1_sb_4__8__chanx_right_out;
wire [0:64] tile_4__9__1_sb_4__8__chany_bottom_out;
wire [0:0] tile_5__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_5__8__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_6__1__0_cbx_6__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_6__1__0_cbx_6__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_6__1__0_cbx_6__0__chanx_left_out;
wire [0:64] tile_6__1__0_cby_6__1__chany_top_out;
wire [0:0] tile_6__1__0_ccff_tail;
wire [0:0] tile_6__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_6__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_6__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_6__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_6__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_6__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_6__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_6__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_6__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_6__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_6__1__0_sb_6__0__chanx_right_out;
wire [0:0] tile_6__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_6__2__0_cbx_6__1__chanx_left_out;
wire [0:64] tile_6__2__0_cby_6__2__chany_top_out;
wire [0:0] tile_6__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_6__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_6__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_6__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_6__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_6__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_6__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_6__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_6__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_6__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_6__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_6__2__0_sb_6__1__chanx_right_out;
wire [0:64] tile_6__2__0_sb_6__1__chany_bottom_out;
wire [0:0] tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_6__2__1_cbx_6__1__chanx_left_out;
wire [0:64] tile_6__2__1_cby_6__2__chany_top_out;
wire [0:0] tile_6__2__1_ccff_tail;
wire [0:0] tile_6__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_6__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_6__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_6__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_6__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_6__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_6__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_6__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_6__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_6__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_6__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_6__2__1_sb_6__1__chanx_right_out;
wire [0:64] tile_6__2__1_sb_6__1__chany_bottom_out;
wire [0:0] tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_6__2__2_cbx_6__1__chanx_left_out;
wire [0:64] tile_6__2__2_cby_6__2__chany_top_out;
wire [0:0] tile_6__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_6__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_6__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_6__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_6__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_6__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_6__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_6__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_6__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_6__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_6__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_6__2__2_sb_6__1__chanx_right_out;
wire [0:64] tile_6__2__2_sb_6__1__chany_bottom_out;
wire [0:0] tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_6__2__3_cbx_6__1__chanx_left_out;
wire [0:64] tile_6__2__3_cby_6__2__chany_top_out;
wire [0:0] tile_6__2__3_ccff_tail;
wire [0:0] tile_6__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_6__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_6__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_6__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_6__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_6__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_6__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_6__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_6__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_6__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_6__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_6__2__3_sb_6__1__chanx_right_out;
wire [0:64] tile_6__2__3_sb_6__1__chany_bottom_out;
wire [0:0] tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_6__2__4_cbx_6__1__chanx_left_out;
wire [0:64] tile_6__2__4_cby_6__2__chany_top_out;
wire [0:0] tile_6__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_6__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_6__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_6__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_6__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_6__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_6__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_6__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_6__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_6__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_6__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_6__2__4_sb_6__1__chanx_right_out;
wire [0:64] tile_6__2__4_sb_6__1__chany_bottom_out;
wire [0:0] tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_6__2__5_cbx_6__1__chanx_left_out;
wire [0:64] tile_6__2__5_cby_6__2__chany_top_out;
wire [0:0] tile_6__2__5_ccff_tail;
wire [0:0] tile_6__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_6__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_6__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_6__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_6__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_6__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_6__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_6__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_6__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_6__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_6__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_6__2__5_sb_6__1__chanx_right_out;
wire [0:64] tile_6__2__5_sb_6__1__chany_bottom_out;
wire [0:0] tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_6__2__6_cbx_6__1__chanx_left_out;
wire [0:64] tile_6__2__6_cby_6__2__chany_top_out;
wire [0:0] tile_6__2__6_ccff_tail;
wire [0:0] tile_6__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] tile_6__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] tile_6__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] tile_6__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] tile_6__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] tile_6__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] tile_6__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] tile_6__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] tile_6__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] tile_6__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] tile_6__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_;
wire [0:64] tile_6__2__6_sb_6__1__chanx_right_out;
wire [0:64] tile_6__2__6_sb_6__1__chany_bottom_out;
wire [0:0] tile_6__8__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
wire [0:0] tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
wire [0:0] tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
wire [0:0] tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
wire [0:0] tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
wire [0:0] tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
wire [0:0] tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
wire [0:0] tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
wire [0:0] tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
wire [0:0] tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
wire [0:0] tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
wire [0:0] tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
wire [0:64] tile_6__9__0_cbx_6__8__chanx_left_out;
wire [0:0] tile_6__9__0_ccff_tail;
wire [0:0] tile_6__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_6__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_6__9__0_sb_6__8__chanx_right_out;
wire [0:64] tile_6__9__0_sb_6__8__chany_bottom_out;
wire [0:0] tile_7__1__0_cbx_7__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_7__1__0_cbx_7__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_7__1__0_cbx_7__0__chanx_left_out;
wire [0:0] tile_7__1__0_cbx_8__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_7__1__0_cbx_8__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:64] tile_7__1__0_cby_8__1__chany_top_out;
wire [0:0] tile_7__1__0_cby_8__1__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_7__1__0_cby_8__1__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:0] tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_7__2__0_cbx_7__1__chanx_left_out;
wire [0:64] tile_7__2__0_cby_8__2__chany_top_out;
wire [0:0] tile_7__2__0_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_7__2__0_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_7__2__0_ccff_tail;
wire [0:0] tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_7__2__0_sb_8__1__chany_bottom_out;
wire [0:0] tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_7__2__1_cbx_7__1__chanx_left_out;
wire [0:64] tile_7__2__1_cby_8__2__chany_top_out;
wire [0:0] tile_7__2__1_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_7__2__1_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_7__2__1_sb_8__1__chany_bottom_out;
wire [0:0] tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_7__2__2_cbx_7__1__chanx_left_out;
wire [0:64] tile_7__2__2_cby_8__2__chany_top_out;
wire [0:0] tile_7__2__2_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_7__2__2_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_7__2__2_ccff_tail;
wire [0:0] tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_7__2__2_sb_8__1__chany_bottom_out;
wire [0:0] tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_7__2__3_cbx_7__1__chanx_left_out;
wire [0:64] tile_7__2__3_cby_8__2__chany_top_out;
wire [0:0] tile_7__2__3_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_7__2__3_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_7__2__3_sb_8__1__chany_bottom_out;
wire [0:0] tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_7__2__4_cbx_7__1__chanx_left_out;
wire [0:64] tile_7__2__4_cby_8__2__chany_top_out;
wire [0:0] tile_7__2__4_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_7__2__4_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_7__2__4_ccff_tail;
wire [0:0] tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_7__2__4_sb_8__1__chany_bottom_out;
wire [0:0] tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_7__2__5_cbx_7__1__chanx_left_out;
wire [0:64] tile_7__2__5_cby_8__2__chany_top_out;
wire [0:0] tile_7__2__5_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_7__2__5_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_7__2__5_sb_8__1__chany_bottom_out;
wire [0:0] tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_7__2__6_cbx_7__1__chanx_left_out;
wire [0:64] tile_7__2__6_cby_8__2__chany_top_out;
wire [0:0] tile_7__2__6_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] tile_7__2__6_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] tile_7__2__6_ccff_tail;
wire [0:0] tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_;
wire [0:0] tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_;
wire [0:0] tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_;
wire [0:0] tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_;
wire [0:0] tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_;
wire [0:0] tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_;
wire [0:0] tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_;
wire [0:0] tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_;
wire [0:64] tile_7__2__6_sb_8__1__chany_bottom_out;
wire [0:0] tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_;
wire [0:0] tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_;
wire [0:0] tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_;
wire [0:0] tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_;
wire [0:0] tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_;
wire [0:0] tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_;
wire [0:0] tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_;
wire [0:0] tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_;
wire [0:64] tile_7__9__0_cbx_7__8__chanx_left_out;
wire [0:0] tile_7__9__0_ccff_tail;
wire [0:0] tile_7__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_7__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_7__9__0_sb_7__8__chanx_right_out;
wire [0:64] tile_8__9__0_cbx_8__8__chanx_left_out;
wire [0:0] tile_8__9__0_ccff_tail;
wire [0:0] tile_8__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_8__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:64] tile_8__9__0_sb_8__8__chany_bottom_out;
wire [0:0] tile_9__1__0_ccff_tail;
wire [0:0] tile_9__1__0_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_9__1__0_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_9__1__1_ccff_tail;
wire [0:0] tile_9__1__1_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_9__1__1_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_9__1__2_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_9__1__2_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_9__1__3_ccff_tail;
wire [0:0] tile_9__1__3_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_9__1__3_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_9__1__4_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_9__1__4_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_9__1__5_ccff_tail;
wire [0:0] tile_9__1__5_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_9__1__5_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_9__1__6_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_9__1__6_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] tile_9__1__7_ccff_tail;
wire [0:0] tile_9__1__7_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] tile_9__1__7_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	tile_0__9_ tile_0__9_ (
		.prog_clk(prog_clk),
		.sb_0__8__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__8__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__8__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__6_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__8__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__6_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__8__chanx_right_in(tile_1__9__0_cbx_1__8__chanx_left_out[0:64]),
		.sb_0__8__chany_bottom_in(tile_0__2__6_cby_0__2__chany_top_out[0:64]),
		.ccff_head(tile_1__9__0_ccff_tail),
		.sb_0__8__chanx_right_out(tile_0__9__0_sb_0__8__chanx_right_out[0:64]),
		.sb_0__8__chany_bottom_out(tile_0__9__0_sb_0__8__chany_bottom_out[0:64]),
		.ccff_tail(ccff_tail[31]));

	tile_1__9_ tile_1__9_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[0:1]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[0:1]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[0:1]),
		.sb_1__8__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_2__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__8__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_2__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__8__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__8__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__8__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__8__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__8__chanx_right_in(tile_2__9__0_cbx_2__8__chanx_left_out[0:64]),
		.sb_1__8__chany_bottom_in(tile_1__2__6_cby_1__2__chany_top_out[0:64]),
		.cbx_1__8__chanx_left_in(tile_0__9__0_sb_0__8__chanx_right_out[0:64]),
		.ccff_head(tile_2__9__0_ccff_tail),
		.cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__8__chanx_right_out(tile_1__9__0_sb_1__8__chanx_right_out[0:64]),
		.sb_1__8__chany_bottom_out(tile_1__9__0_sb_1__8__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_1__8__chanx_left_out(tile_1__9__0_cbx_1__8__chanx_left_out[0:64]),
		.ccff_tail(tile_1__9__0_ccff_tail));

	tile_2__9_ tile_2__9_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[2:3]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[2:3]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[2:3]),
		.sb_2__8__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_3__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_2__8__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_3__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_2__8__chanx_right_in(tile_3__9__0_cbx_3__8__chanx_left_out[0:64]),
		.cbx_2__8__chanx_left_in(tile_1__9__0_sb_1__8__chanx_right_out[0:64]),
		.ccff_head(tile_3__9__0_ccff_tail),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.sb_2__8__chanx_right_out(tile_2__9__0_sb_2__8__chanx_right_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_2__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_2__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_2__8__chanx_left_out(tile_2__9__0_cbx_2__8__chanx_left_out[0:64]),
		.ccff_tail(tile_2__9__0_ccff_tail));

	tile_3__9_ tile_3__9_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[4:5]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[4:5]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[4:5]),
		.sb_3__8__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_4__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_3__8__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_4__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_3__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_3__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_3__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_3__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_3__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_3__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_3__8__chanx_right_in(tile_4__9__0_cbx_4__8__chanx_left_out[0:64]),
		.sb_3__8__chany_bottom_in(tile_2__2__6_cby_3__2__chany_top_out[0:64]),
		.cbx_3__8__chanx_left_in(tile_2__9__0_sb_2__8__chanx_right_out[0:64]),
		.ccff_head(tile_4__9__0_ccff_tail),
		.sb_3__8__chanx_right_out(tile_3__9__0_sb_3__8__chanx_right_out[0:64]),
		.sb_3__8__chany_bottom_out(tile_3__9__0_sb_3__8__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_3__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_3__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_3__8__chanx_left_out(tile_3__9__0_cbx_3__8__chanx_left_out[0:64]),
		.ccff_tail(tile_3__9__0_ccff_tail));

	tile_4__9_ tile_4__9_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[6:7]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[6:7]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[6:7]),
		.sb_4__8__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_4__9__1_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_4__8__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_4__9__1_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_4__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__8__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_4__8__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_4__8__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_4__8__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_4__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__8__chanx_right_in(tile_4__9__1_cbx_4__8__chanx_left_out[0:64]),
		.sb_4__8__chany_bottom_in(tile_4__2__6_cby_4__2__chany_top_out[0:64]),
		.cbx_4__8__chanx_left_in(tile_3__9__0_sb_3__8__chanx_right_out[0:64]),
		.ccff_head(tile_4__9__1_ccff_tail),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_4__8__chanx_right_out(tile_4__9__0_sb_4__8__chanx_right_out[0:64]),
		.sb_4__8__chany_bottom_out(tile_4__9__0_sb_4__8__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_4__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_4__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_4__8__chanx_left_out(tile_4__9__0_cbx_4__8__chanx_left_out[0:64]),
		.ccff_tail(tile_4__9__0_ccff_tail));

	tile_4__9_ tile_5__9_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[8:9]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[8:9]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[8:9]),
		.sb_4__8__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_6__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_4__8__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_6__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_4__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__8__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_4__8__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_4__8__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_4__8__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_4__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__8__chanx_right_in(tile_6__9__0_cbx_6__8__chanx_left_out[0:64]),
		.sb_4__8__chany_bottom_in(tile_4__2__13_cby_4__2__chany_top_out[0:64]),
		.cbx_4__8__chanx_left_in(tile_4__9__0_sb_4__8__chanx_right_out[0:64]),
		.ccff_head(tile_6__9__0_ccff_tail),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_4__8__chanx_right_out(tile_4__9__1_sb_4__8__chanx_right_out[0:64]),
		.sb_4__8__chany_bottom_out(tile_4__9__1_sb_4__8__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_4__9__1_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_4__9__1_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_4__8__chanx_left_out(tile_4__9__1_cbx_4__8__chanx_left_out[0:64]),
		.ccff_tail(tile_4__9__1_ccff_tail));

	tile_6__9_ tile_6__9_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[10:11]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[10:11]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[10:11]),
		.sb_6__8__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_7__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_6__8__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_7__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_6__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_6__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_6__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_6__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_6__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_6__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_6__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_6__8__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_6__8__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_6__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_6__8__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_6__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_6__8__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_6__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_6__8__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_6__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_6__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_6__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_6__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_6__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_6__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_6__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_6__8__chanx_right_in(tile_7__9__0_cbx_7__8__chanx_left_out[0:64]),
		.sb_6__8__chany_bottom_in(tile_6__2__6_cby_6__2__chany_top_out[0:64]),
		.cbx_6__8__chanx_left_in(tile_4__9__1_sb_4__8__chanx_right_out[0:64]),
		.ccff_head(tile_7__9__0_ccff_tail),
		.cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_6__8__chanx_right_out(tile_6__9__0_sb_6__8__chanx_right_out[0:64]),
		.sb_6__8__chany_bottom_out(tile_6__9__0_sb_6__8__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_6__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_6__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_6__8__chanx_left_out(tile_6__9__0_cbx_6__8__chanx_left_out[0:64]),
		.ccff_tail(tile_6__9__0_ccff_tail));

	tile_7__9_ tile_7__9_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[12:13]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[12:13]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[12:13]),
		.sb_7__8__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_8__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_7__8__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_8__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_7__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_7__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_7__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_7__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_7__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_7__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_7__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_7__8__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_7__8__chanx_right_in(tile_8__9__0_cbx_8__8__chanx_left_out[0:64]),
		.cbx_7__8__chanx_left_in(tile_6__9__0_sb_6__8__chanx_right_out[0:64]),
		.ccff_head(tile_8__9__0_ccff_tail),
		.cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.sb_7__8__chanx_right_out(tile_7__9__0_sb_7__8__chanx_right_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_7__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_7__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_7__8__chanx_left_out(tile_7__9__0_cbx_7__8__chanx_left_out[0:64]),
		.ccff_tail(tile_7__9__0_ccff_tail));

	tile_8__9_ tile_8__9_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[14:15]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[14:15]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[14:15]),
		.sb_8__8__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__0_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_8__8__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__0_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_8__8__chany_bottom_in(tile_7__2__6_cby_8__2__chany_top_out[0:64]),
		.cbx_8__8__chanx_left_in(tile_7__9__0_sb_7__8__chanx_right_out[0:64]),
		.ccff_head(tile_9__1__0_ccff_tail),
		.sb_8__8__chany_bottom_out(tile_8__9__0_sb_8__8__chany_bottom_out[0:64]),
		.grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_8__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_8__9__0_grid_io_top_top_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.cbx_8__8__chanx_left_out(tile_8__9__0_cbx_8__8__chanx_left_out[0:64]),
		.ccff_tail(tile_8__9__0_ccff_tail));

	tile_9__1_ tile_9__8_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[16:17]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[16:17]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[16:17]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__2__6_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__2__6_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_7__2__6_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__0_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__0_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_9__1__0_ccff_tail));

	tile_9__1_ tile_9__7_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[18:19]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[18:19]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[18:19]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__2__5_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__2__5_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(ccff_head[28]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__1_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__1_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_9__1__1_ccff_tail));

	tile_9__1_ tile_9__6_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[20:21]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[20:21]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[20:21]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__2__4_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__2__4_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_7__2__4_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__2_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__2_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(ccff_tail[27]));

	tile_9__1_ tile_9__5_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[22:23]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[22:23]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[22:23]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__2__3_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__2__3_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(ccff_head[20]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__3_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__3_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_9__1__3_ccff_tail));

	tile_9__1_ tile_9__4_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[24:25]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[24:25]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[24:25]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__2__2_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__2__2_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_7__2__2_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__4_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__4_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(ccff_tail[19]));

	tile_9__1_ tile_9__3_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[26:27]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[26:27]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[26:27]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__2__1_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__2__1_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(ccff_head[12]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__5_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__5_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_9__1__5_ccff_tail));

	tile_9__1_ tile_9__2_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[28:29]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[28:29]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[28:29]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__2__0_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__2__0_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_7__2__0_ccff_tail),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__6_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__6_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(ccff_tail[11]));

	tile_9__1_ tile_9__1_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[30:31]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[30:31]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[30:31]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__1__0_cby_8__1__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__1__0_cby_8__1__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(ccff_head[4]),
		.grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__7_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__7_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_9__1__7_ccff_tail));

	tile_1__0_ tile_8__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[32:33]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[32:33]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[32:33]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__1__0_cbx_8__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__1__0_cbx_8__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__1_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__0_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__0_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(ccff_tail[3]));

	tile_1__0_ tile_7__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[34:35]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[34:35]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[34:35]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__1__0_cbx_7__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__1__0_cbx_7__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(ccff_head[3]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__1_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__1_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__1_ccff_tail));

	tile_1__0_ tile_6__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[36:37]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[36:37]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[36:37]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_6__1__0_cbx_6__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_6__1__0_cbx_6__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__3_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__2_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__2_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(ccff_tail[2]));

	tile_1__0_ tile_5__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[38:39]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[38:39]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[38:39]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_4__1__1_cbx_4__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_4__1__1_cbx_4__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(ccff_head[2]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__3_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__3_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__3_ccff_tail));

	tile_1__0_ tile_4__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[40:41]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[40:41]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[40:41]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_4__1__0_cbx_4__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_4__1__0_cbx_4__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__5_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__4_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__4_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(ccff_tail[1]));

	tile_1__0_ tile_3__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[42:43]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[42:43]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[42:43]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_2__1__0_cbx_3__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_2__1__0_cbx_3__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(ccff_head[1]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__5_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__5_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__5_ccff_tail));

	tile_1__0_ tile_2__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[44:45]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[44:45]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[44:45]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_2__1__0_cbx_2__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_2__1__0_cbx_2__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(tile_1__0__7_ccff_tail),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__6_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__6_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(ccff_tail[0]));

	tile_1__0_ tile_1__0_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[46:47]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[46:47]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[46:47]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__0_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__0_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(ccff_head[0]),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__7_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__7_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.ccff_tail(tile_1__0__7_ccff_tail));

	tile_0__1_ tile_0__1_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[48:49]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[48:49]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[48:49]),
		.sb_0__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__7_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__7_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__0__chanx_right_in(tile_1__1__0_cbx_1__0__chanx_left_out[0:64]),
		.cby_0__1__chany_top_in(tile_0__2__0_sb_0__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__1__0_ccff_tail),
		.sb_0__0__chanx_right_out(tile_0__1__0_sb_0__0__chanx_right_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__1__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__1__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__1__chany_top_out(tile_0__1__0_cby_0__1__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[7]));

	tile_0__2_ tile_0__2_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[50:51]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[50:51]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[50:51]),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__1__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__1__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__1__chanx_right_in(tile_1__2__0_cbx_1__1__chanx_left_out[0:64]),
		.sb_0__1__chany_bottom_in(tile_0__1__0_cby_0__1__chany_top_out[0:64]),
		.cby_0__2__chany_top_in(tile_0__2__1_sb_0__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[8]),
		.sb_0__1__chanx_right_out(tile_0__2__0_sb_0__1__chanx_right_out[0:64]),
		.sb_0__1__chany_bottom_out(tile_0__2__0_sb_0__1__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__2__chany_top_out(tile_0__2__0_cby_0__2__chany_top_out[0:64]),
		.ccff_tail(tile_0__2__0_ccff_tail));

	tile_0__2_ tile_0__3_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[52:53]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[52:53]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[52:53]),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__0_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__0_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__1__chanx_right_in(tile_1__2__1_cbx_1__1__chanx_left_out[0:64]),
		.sb_0__1__chany_bottom_in(tile_0__2__0_cby_0__2__chany_top_out[0:64]),
		.cby_0__2__chany_top_in(tile_0__2__2_sb_0__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__1_ccff_tail),
		.sb_0__1__chanx_right_out(tile_0__2__1_sb_0__1__chanx_right_out[0:64]),
		.sb_0__1__chany_bottom_out(tile_0__2__1_sb_0__1__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__1_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__1_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__2__chany_top_out(tile_0__2__1_cby_0__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[15]));

	tile_0__2_ tile_0__4_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[54:55]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[54:55]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[54:55]),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__1_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__1_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__1__chanx_right_in(tile_1__2__2_cbx_1__1__chanx_left_out[0:64]),
		.sb_0__1__chany_bottom_in(tile_0__2__1_cby_0__2__chany_top_out[0:64]),
		.cby_0__2__chany_top_in(tile_0__2__3_sb_0__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[16]),
		.sb_0__1__chanx_right_out(tile_0__2__2_sb_0__1__chanx_right_out[0:64]),
		.sb_0__1__chany_bottom_out(tile_0__2__2_sb_0__1__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__2_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__2_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__2__chany_top_out(tile_0__2__2_cby_0__2__chany_top_out[0:64]),
		.ccff_tail(tile_0__2__2_ccff_tail));

	tile_0__2_ tile_0__5_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[56:57]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[56:57]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[56:57]),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__2_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__2_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__1__chanx_right_in(tile_1__2__3_cbx_1__1__chanx_left_out[0:64]),
		.sb_0__1__chany_bottom_in(tile_0__2__2_cby_0__2__chany_top_out[0:64]),
		.cby_0__2__chany_top_in(tile_0__2__4_sb_0__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__3_ccff_tail),
		.sb_0__1__chanx_right_out(tile_0__2__3_sb_0__1__chanx_right_out[0:64]),
		.sb_0__1__chany_bottom_out(tile_0__2__3_sb_0__1__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__3_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__3_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__2__chany_top_out(tile_0__2__3_cby_0__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[23]));

	tile_0__2_ tile_0__6_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[58:59]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[58:59]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[58:59]),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__3_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__3_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__1__chanx_right_in(tile_1__2__4_cbx_1__1__chanx_left_out[0:64]),
		.sb_0__1__chany_bottom_in(tile_0__2__3_cby_0__2__chany_top_out[0:64]),
		.cby_0__2__chany_top_in(tile_0__2__5_sb_0__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[24]),
		.sb_0__1__chanx_right_out(tile_0__2__4_sb_0__1__chanx_right_out[0:64]),
		.sb_0__1__chany_bottom_out(tile_0__2__4_sb_0__1__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__4_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__4_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__2__chany_top_out(tile_0__2__4_cby_0__2__chany_top_out[0:64]),
		.ccff_tail(tile_0__2__4_ccff_tail));

	tile_0__2_ tile_0__7_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[60:61]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[60:61]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[60:61]),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__4_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__4_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__1__chanx_right_in(tile_1__2__5_cbx_1__1__chanx_left_out[0:64]),
		.sb_0__1__chany_bottom_in(tile_0__2__4_cby_0__2__chany_top_out[0:64]),
		.cby_0__2__chany_top_in(tile_0__2__6_sb_0__1__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__5_ccff_tail),
		.sb_0__1__chanx_right_out(tile_0__2__5_sb_0__1__chanx_right_out[0:64]),
		.sb_0__1__chany_bottom_out(tile_0__2__5_sb_0__1__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__5_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__5_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__2__chany_top_out(tile_0__2__5_cby_0__2__chany_top_out[0:64]),
		.ccff_tail(tile_0__2__5_ccff_tail));

	tile_0__2_ tile_0__8_ (
		.IO_ISOL_N(IO_ISOL_N),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[62:63]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[62:63]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[62:63]),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__5_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_0__1__bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__5_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_0__1__chanx_right_in(tile_1__2__6_cbx_1__1__chanx_left_out[0:64]),
		.sb_0__1__chany_bottom_in(tile_0__2__5_cby_0__2__chany_top_out[0:64]),
		.cby_0__2__chany_top_in(tile_0__9__0_sb_0__8__chany_bottom_out[0:64]),
		.ccff_head(tile_0__2__5_ccff_tail),
		.sb_0__1__chanx_right_out(tile_0__2__6_sb_0__1__chanx_right_out[0:64]),
		.sb_0__1__chany_bottom_out(tile_0__2__6_sb_0__1__chany_bottom_out[0:64]),
		.grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_(tile_0__2__6_grid_io_left_left_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_(tile_0__2__6_grid_io_left_left_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.cby_0__2__chany_top_out(tile_0__2__6_cby_0__2__chany_top_out[0:64]),
		.ccff_tail(tile_0__2__6_ccff_tail));

	tile_1__1_ tile_1__1_ (
		.prog_clk(prog_clk),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.sb_1__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__6_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__6_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__7_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_1__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__7_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_1__0__chanx_right_in(tile_2__1__0_cbx_2__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_0_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_1__0__chanx_left_in(tile_0__1__0_sb_0__0__chanx_right_out[0:64]),
		.cby_1__1__chany_top_in(tile_1__2__0_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[7]),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_1__1__0_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_1__1__0_cbx_1__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_1__0__chanx_right_out(tile_1__1__0_sb_1__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__0__chanx_left_out(tile_1__1__0_cbx_1__0__chanx_left_out[0:64]),
		.cby_1__1__chany_top_out(tile_1__1__0_cby_1__1__chany_top_out[0:64]),
		.ccff_tail(tile_1__1__0_ccff_tail));

	tile_1__2_ tile_1__2_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_2__2__0_cbx_2__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__1__0_cby_1__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_1_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_1__1__chanx_left_in(tile_0__2__0_sb_0__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__1_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_0__2__0_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__0_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__0_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__0_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__0_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__0_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[8]));

	tile_1__2_ tile_1__3_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_2__2__1_cbx_2__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__0_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_2_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_1__1__chanx_left_in(tile_0__2__1_sb_0__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__2_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[15]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__1_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__1_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__1_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__1_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__1_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__1_ccff_tail));

	tile_1__2_ tile_1__4_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_2__2__2_cbx_2__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__1_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_3_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_1__1__chanx_left_in(tile_0__2__2_sb_0__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__3_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_0__2__2_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__2_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__2_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__2_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__2_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__2_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[16]));

	tile_1__2_ tile_1__5_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_2__2__3_cbx_2__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__2_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_4_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_1__1__chanx_left_in(tile_0__2__3_sb_0__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__4_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[23]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__3_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__3_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__3_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__3_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__3_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__3_ccff_tail));

	tile_1__2_ tile_1__6_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_2__2__4_cbx_2__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__3_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_5_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_1__1__chanx_left_in(tile_0__2__4_sb_0__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__5_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(tile_0__2__4_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__4_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__4_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__4_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__4_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__4_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[24]));

	tile_1__2_ tile_1__7_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_2__2__5_cbx_2__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__4_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_6_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_1__1__chanx_left_in(tile_0__2__5_sb_0__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__2__6_sb_1__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[31]),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__5_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__5_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__5_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__5_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__5_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__5_ccff_tail));

	tile_1__2_ tile_1__8_ (
		.prog_clk(prog_clk),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.sb_1__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_1__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_1__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_1__1__chanx_right_in(tile_2__2__6_cbx_2__1__chanx_left_out[0:64]),
		.sb_1__1__chany_bottom_in(tile_1__2__5_cby_1__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__9__0_cbx_1__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_1__8__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_1__1__chanx_left_in(tile_0__2__6_sb_0__1__chanx_right_out[0:64]),
		.cby_1__2__chany_top_in(tile_1__9__0_sb_1__8__chany_bottom_out[0:64]),
		.ccff_head(tile_0__2__6_ccff_tail),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_1__2__6_cbx_1__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_1__1__chanx_right_out(tile_1__2__6_sb_1__1__chanx_right_out[0:64]),
		.sb_1__1__chany_bottom_out(tile_1__2__6_sb_1__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_1__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_1__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_1__1__chanx_left_out(tile_1__2__6_cbx_1__1__chanx_left_out[0:64]),
		.cby_1__2__chany_top_out(tile_1__2__6_cby_1__2__chany_top_out[0:64]),
		.ccff_tail(tile_1__2__6_ccff_tail));

	tile_2__1_ tile_2__1_ (
		.prog_clk(prog_clk),
		.sb_2__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__5_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_2__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__5_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_2__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__6_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_2__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__6_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_3__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_3__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_3__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_3__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_3__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_3__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_3__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__4_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_3__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__4_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_3__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__5_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_3__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__5_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_3__0__chanx_right_in(tile_4__1__0_cbx_4__0__chanx_left_out[0:64]),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.cbx_2__0__chanx_left_in(tile_1__1__0_sb_1__0__chanx_right_out[0:64]),
		.cby_3__1__chany_top_in(tile_2__2__0_sb_3__1__chany_bottom_out[0:64]),
		.ccff_head(tile_4__1__0_ccff_tail),
		.cbx_2__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_2__1__0_cbx_2__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_2__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_2__1__0_cbx_2__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.cbx_3__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_2__1__0_cbx_3__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_3__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_2__1__0_cbx_3__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_3__0__chanx_right_out(tile_2__1__0_sb_3__0__chanx_right_out[0:64]),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_2__1__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.cbx_2__0__chanx_left_out(tile_2__1__0_cbx_2__0__chanx_left_out[0:64]),
		.cby_3__1__chany_top_out(tile_2__1__0_cby_3__1__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[6]));

	tile_2__2_ tile_2__2_ (
		.prog_clk(prog_clk),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_3__1__chanx_right_in(tile_4__2__0_cbx_4__1__chanx_left_out[0:64]),
		.sb_3__1__chany_bottom_in(tile_2__1__0_cby_3__1__chany_top_out[0:64]),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.cbx_2__1__chanx_left_in(tile_1__2__0_sb_1__1__chanx_right_out[0:64]),
		.cby_3__2__chany_top_in(tile_2__2__1_sb_3__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[9]),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_(tile_2__2__0_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.sb_3__1__chanx_right_out(tile_2__2__0_sb_3__1__chanx_right_out[0:64]),
		.sb_3__1__chany_bottom_out(tile_2__2__0_sb_3__1__chany_bottom_out[0:64]),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_2__2__0_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.cbx_2__1__chanx_left_out(tile_2__2__0_cbx_2__1__chanx_left_out[0:64]),
		.cby_3__2__chany_top_out(tile_2__2__0_cby_3__2__chany_top_out[0:64]),
		.ccff_tail(tile_2__2__0_ccff_tail));

	tile_2__2_ tile_2__3_ (
		.prog_clk(prog_clk),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_3__1__chanx_right_in(tile_4__2__1_cbx_4__1__chanx_left_out[0:64]),
		.sb_3__1__chany_bottom_in(tile_2__2__0_cby_3__2__chany_top_out[0:64]),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.cbx_2__1__chanx_left_in(tile_1__2__1_sb_1__1__chanx_right_out[0:64]),
		.cby_3__2__chany_top_in(tile_2__2__2_sb_3__1__chany_bottom_out[0:64]),
		.ccff_head(tile_4__2__1_ccff_tail),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_(tile_2__2__1_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.sb_3__1__chanx_right_out(tile_2__2__1_sb_3__1__chanx_right_out[0:64]),
		.sb_3__1__chany_bottom_out(tile_2__2__1_sb_3__1__chany_bottom_out[0:64]),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_2__2__1_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.cbx_2__1__chanx_left_out(tile_2__2__1_cbx_2__1__chanx_left_out[0:64]),
		.cby_3__2__chany_top_out(tile_2__2__1_cby_3__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[14]));

	tile_2__2_ tile_2__4_ (
		.prog_clk(prog_clk),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_3__1__chanx_right_in(tile_4__2__2_cbx_4__1__chanx_left_out[0:64]),
		.sb_3__1__chany_bottom_in(tile_2__2__1_cby_3__2__chany_top_out[0:64]),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.cbx_2__1__chanx_left_in(tile_1__2__2_sb_1__1__chanx_right_out[0:64]),
		.cby_3__2__chany_top_in(tile_2__2__3_sb_3__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[17]),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_(tile_2__2__2_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.sb_3__1__chanx_right_out(tile_2__2__2_sb_3__1__chanx_right_out[0:64]),
		.sb_3__1__chany_bottom_out(tile_2__2__2_sb_3__1__chany_bottom_out[0:64]),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_2__2__2_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.cbx_2__1__chanx_left_out(tile_2__2__2_cbx_2__1__chanx_left_out[0:64]),
		.cby_3__2__chany_top_out(tile_2__2__2_cby_3__2__chany_top_out[0:64]),
		.ccff_tail(tile_2__2__2_ccff_tail));

	tile_2__2_ tile_2__5_ (
		.prog_clk(prog_clk),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_3__1__chanx_right_in(tile_4__2__3_cbx_4__1__chanx_left_out[0:64]),
		.sb_3__1__chany_bottom_in(tile_2__2__2_cby_3__2__chany_top_out[0:64]),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.cbx_2__1__chanx_left_in(tile_1__2__3_sb_1__1__chanx_right_out[0:64]),
		.cby_3__2__chany_top_in(tile_2__2__4_sb_3__1__chany_bottom_out[0:64]),
		.ccff_head(tile_4__2__3_ccff_tail),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_(tile_2__2__3_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.sb_3__1__chanx_right_out(tile_2__2__3_sb_3__1__chanx_right_out[0:64]),
		.sb_3__1__chany_bottom_out(tile_2__2__3_sb_3__1__chany_bottom_out[0:64]),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_2__2__3_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.cbx_2__1__chanx_left_out(tile_2__2__3_cbx_2__1__chanx_left_out[0:64]),
		.cby_3__2__chany_top_out(tile_2__2__3_cby_3__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[22]));

	tile_2__2_ tile_2__6_ (
		.prog_clk(prog_clk),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_3__1__chanx_right_in(tile_4__2__4_cbx_4__1__chanx_left_out[0:64]),
		.sb_3__1__chany_bottom_in(tile_2__2__3_cby_3__2__chany_top_out[0:64]),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.cbx_2__1__chanx_left_in(tile_1__2__4_sb_1__1__chanx_right_out[0:64]),
		.cby_3__2__chany_top_in(tile_2__2__5_sb_3__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[25]),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_(tile_2__2__4_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.sb_3__1__chanx_right_out(tile_2__2__4_sb_3__1__chanx_right_out[0:64]),
		.sb_3__1__chany_bottom_out(tile_2__2__4_sb_3__1__chany_bottom_out[0:64]),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_2__2__4_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.cbx_2__1__chanx_left_out(tile_2__2__4_cbx_2__1__chanx_left_out[0:64]),
		.cby_3__2__chany_top_out(tile_2__2__4_cby_3__2__chany_top_out[0:64]),
		.ccff_tail(tile_2__2__4_ccff_tail));

	tile_2__2_ tile_2__7_ (
		.prog_clk(prog_clk),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_3__1__chanx_right_in(tile_4__2__5_cbx_4__1__chanx_left_out[0:64]),
		.sb_3__1__chany_bottom_in(tile_2__2__4_cby_3__2__chany_top_out[0:64]),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.cbx_2__1__chanx_left_in(tile_1__2__5_sb_1__1__chanx_right_out[0:64]),
		.cby_3__2__chany_top_in(tile_2__2__6_sb_3__1__chany_bottom_out[0:64]),
		.ccff_head(tile_4__2__5_ccff_tail),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_(tile_2__2__5_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.sb_3__1__chanx_right_out(tile_2__2__5_sb_3__1__chanx_right_out[0:64]),
		.sb_3__1__chany_bottom_out(tile_2__2__5_sb_3__1__chany_bottom_out[0:64]),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_2__2__5_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.cbx_2__1__chanx_left_out(tile_2__2__5_cbx_2__1__chanx_left_out[0:64]),
		.cby_3__2__chany_top_out(tile_2__2__5_cby_3__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[30]));

	tile_2__2_ tile_2__8_ (
		.prog_clk(prog_clk),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_3__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_3__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_3__1__chanx_right_in(tile_4__2__6_cbx_4__1__chanx_left_out[0:64]),
		.sb_3__1__chany_bottom_in(tile_2__2__5_cby_3__2__chany_top_out[0:64]),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_(tile_2__9__0_cbx_2__8__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.cbx_2__1__chanx_left_in(tile_1__2__6_sb_1__1__chanx_right_out[0:64]),
		.cby_3__2__chany_top_in(tile_3__9__0_sb_3__8__chany_bottom_out[0:64]),
		.ccff_head(tile_1__2__6_ccff_tail),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_sign_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_1_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_2_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_3_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_4_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_5_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_6_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_7_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_8_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_9_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_10_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_11_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_12_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_13_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_14_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_15_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_16_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_17_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_a_18_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_0_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_1_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_2_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_3_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_4_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_5_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_6_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_7_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_8_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_9_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_10_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_11_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_12_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_13_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_14_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_15_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_16_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_17_),
		.cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_(tile_2__2__6_cbx_2__1__bottom_grid_top_width_0_height_0_subtile_0__pin_b_18_),
		.sb_3__1__chanx_right_out(tile_2__2__6_sb_3__1__chanx_right_out[0:64]),
		.sb_3__1__chany_bottom_out(tile_2__2__6_sb_3__1__chany_bottom_out[0:64]),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_(tile_2__2__6_grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.cbx_2__1__chanx_left_out(tile_2__2__6_cbx_2__1__chanx_left_out[0:64]),
		.cby_3__2__chany_top_out(tile_2__2__6_cby_3__2__chany_top_out[0:64]),
		.ccff_tail(tile_2__2__6_ccff_tail));

	tile_4__1_ tile_4__1_ (
		.prog_clk(prog_clk),
		.sb_4__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_4__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_4__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_4__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_4__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_4__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_4__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__3_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_4__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__3_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_4__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__4_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_4__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__4_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_4__0__chanx_right_in(tile_4__1__1_cbx_4__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_7_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_4__0__chanx_left_in(tile_2__1__0_sb_3__0__chanx_right_out[0:64]),
		.cby_4__1__chany_top_in(tile_4__2__0_sb_4__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[6]),
		.cbx_4__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_4__1__0_cbx_4__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_4__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_4__1__0_cbx_4__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_4__0__chanx_right_out(tile_4__1__0_sb_4__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_4__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_4__0__chanx_left_out(tile_4__1__0_cbx_4__0__chanx_left_out[0:64]),
		.cby_4__1__chany_top_out(tile_4__1__0_cby_4__1__chany_top_out[0:64]),
		.ccff_tail(tile_4__1__0_ccff_tail));

	tile_4__1_ tile_5__1_ (
		.prog_clk(prog_clk),
		.sb_4__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_6__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_4__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_6__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_4__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_6__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_4__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_6__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_4__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_6__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_4__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_6__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_4__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__2_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_4__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__2_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_4__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__3_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_4__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__3_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_4__0__chanx_right_in(tile_6__1__0_cbx_6__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_14_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_4__0__chanx_left_in(tile_4__1__0_sb_4__0__chanx_right_out[0:64]),
		.cby_4__1__chany_top_in(tile_4__2__7_sb_4__1__chany_bottom_out[0:64]),
		.ccff_head(tile_6__1__0_ccff_tail),
		.cbx_4__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_4__1__1_cbx_4__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_4__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_4__1__1_cbx_4__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_4__0__chanx_right_out(tile_4__1__1_sb_4__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_5__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__1__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_4__0__chanx_left_out(tile_4__1__1_cbx_4__0__chanx_left_out[0:64]),
		.cby_4__1__chany_top_out(tile_4__1__1_cby_4__1__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[5]));

	tile_4__2_ tile_4__2_ (
		.prog_clk(prog_clk),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__chanx_right_in(tile_4__2__7_cbx_4__1__chanx_left_out[0:64]),
		.sb_4__1__chany_bottom_in(tile_4__1__0_cby_4__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_8_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_4__1__chanx_left_in(tile_2__2__0_sb_3__1__chanx_right_out[0:64]),
		.cby_4__2__chany_top_in(tile_4__2__1_sb_4__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__2__0_ccff_tail),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__0_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_4__1__chanx_right_out(tile_4__2__0_sb_4__1__chanx_right_out[0:64]),
		.sb_4__1__chany_bottom_out(tile_4__2__0_sb_4__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_4__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_4__1__chanx_left_out(tile_4__2__0_cbx_4__1__chanx_left_out[0:64]),
		.cby_4__2__chany_top_out(tile_4__2__0_cby_4__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[9]));

	tile_4__2_ tile_4__3_ (
		.prog_clk(prog_clk),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__chanx_right_in(tile_4__2__8_cbx_4__1__chanx_left_out[0:64]),
		.sb_4__1__chany_bottom_in(tile_4__2__0_cby_4__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_9_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_4__1__chanx_left_in(tile_2__2__1_sb_3__1__chanx_right_out[0:64]),
		.cby_4__2__chany_top_in(tile_4__2__2_sb_4__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[14]),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__1_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_4__1__chanx_right_out(tile_4__2__1_sb_4__1__chanx_right_out[0:64]),
		.sb_4__1__chany_bottom_out(tile_4__2__1_sb_4__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_4__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_4__1__chanx_left_out(tile_4__2__1_cbx_4__1__chanx_left_out[0:64]),
		.cby_4__2__chany_top_out(tile_4__2__1_cby_4__2__chany_top_out[0:64]),
		.ccff_tail(tile_4__2__1_ccff_tail));

	tile_4__2_ tile_4__4_ (
		.prog_clk(prog_clk),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__chanx_right_in(tile_4__2__9_cbx_4__1__chanx_left_out[0:64]),
		.sb_4__1__chany_bottom_in(tile_4__2__1_cby_4__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_10_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_4__1__chanx_left_in(tile_2__2__2_sb_3__1__chanx_right_out[0:64]),
		.cby_4__2__chany_top_in(tile_4__2__3_sb_4__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__2__2_ccff_tail),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__2_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_4__1__chanx_right_out(tile_4__2__2_sb_4__1__chanx_right_out[0:64]),
		.sb_4__1__chany_bottom_out(tile_4__2__2_sb_4__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_4__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_4__1__chanx_left_out(tile_4__2__2_cbx_4__1__chanx_left_out[0:64]),
		.cby_4__2__chany_top_out(tile_4__2__2_cby_4__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[17]));

	tile_4__2_ tile_4__5_ (
		.prog_clk(prog_clk),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__chanx_right_in(tile_4__2__10_cbx_4__1__chanx_left_out[0:64]),
		.sb_4__1__chany_bottom_in(tile_4__2__2_cby_4__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_11_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_4__1__chanx_left_in(tile_2__2__3_sb_3__1__chanx_right_out[0:64]),
		.cby_4__2__chany_top_in(tile_4__2__4_sb_4__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[22]),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__3_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_4__1__chanx_right_out(tile_4__2__3_sb_4__1__chanx_right_out[0:64]),
		.sb_4__1__chany_bottom_out(tile_4__2__3_sb_4__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_4__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_4__1__chanx_left_out(tile_4__2__3_cbx_4__1__chanx_left_out[0:64]),
		.cby_4__2__chany_top_out(tile_4__2__3_cby_4__2__chany_top_out[0:64]),
		.ccff_tail(tile_4__2__3_ccff_tail));

	tile_4__2_ tile_4__6_ (
		.prog_clk(prog_clk),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__chanx_right_in(tile_4__2__11_cbx_4__1__chanx_left_out[0:64]),
		.sb_4__1__chany_bottom_in(tile_4__2__3_cby_4__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_12_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_4__1__chanx_left_in(tile_2__2__4_sb_3__1__chanx_right_out[0:64]),
		.cby_4__2__chany_top_in(tile_4__2__5_sb_4__1__chany_bottom_out[0:64]),
		.ccff_head(tile_2__2__4_ccff_tail),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__4_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_4__1__chanx_right_out(tile_4__2__4_sb_4__1__chanx_right_out[0:64]),
		.sb_4__1__chany_bottom_out(tile_4__2__4_sb_4__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_4__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_4__1__chanx_left_out(tile_4__2__4_cbx_4__1__chanx_left_out[0:64]),
		.cby_4__2__chany_top_out(tile_4__2__4_cby_4__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[25]));

	tile_4__2_ tile_4__7_ (
		.prog_clk(prog_clk),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__chanx_right_in(tile_4__2__12_cbx_4__1__chanx_left_out[0:64]),
		.sb_4__1__chany_bottom_in(tile_4__2__4_cby_4__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_13_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_4__1__chanx_left_in(tile_2__2__5_sb_3__1__chanx_right_out[0:64]),
		.cby_4__2__chany_top_in(tile_4__2__6_sb_4__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[30]),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__5_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_4__1__chanx_right_out(tile_4__2__5_sb_4__1__chanx_right_out[0:64]),
		.sb_4__1__chany_bottom_out(tile_4__2__5_sb_4__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_4__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_4__1__chanx_left_out(tile_4__2__5_cbx_4__1__chanx_left_out[0:64]),
		.cby_4__2__chany_top_out(tile_4__2__5_cby_4__2__chany_top_out[0:64]),
		.ccff_tail(tile_4__2__5_ccff_tail));

	tile_4__2_ tile_4__8_ (
		.prog_clk(prog_clk),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__chanx_right_in(tile_4__2__13_cbx_4__1__chanx_left_out[0:64]),
		.sb_4__1__chany_bottom_in(tile_4__2__5_cby_4__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__9__0_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_4__8__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_4__1__chanx_left_in(tile_2__2__6_sb_3__1__chanx_right_out[0:64]),
		.cby_4__2__chany_top_in(tile_4__9__0_sb_4__8__chany_bottom_out[0:64]),
		.ccff_head(tile_2__2__6_ccff_tail),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__6_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_4__1__chanx_right_out(tile_4__2__6_sb_4__1__chanx_right_out[0:64]),
		.sb_4__1__chany_bottom_out(tile_4__2__6_sb_4__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_4__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_4__1__chanx_left_out(tile_4__2__6_cbx_4__1__chanx_left_out[0:64]),
		.cby_4__2__chany_top_out(tile_4__2__6_cby_4__2__chany_top_out[0:64]),
		.ccff_tail(tile_4__2__6_ccff_tail));

	tile_4__2_ tile_5__2_ (
		.prog_clk(prog_clk),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_6__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_6__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_6__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_6__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_6__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_6__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__1__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__1__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__chanx_right_in(tile_6__2__0_cbx_6__1__chanx_left_out[0:64]),
		.sb_4__1__chany_bottom_in(tile_4__1__1_cby_4__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_15_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_4__1__chanx_left_in(tile_4__2__0_sb_4__1__chanx_right_out[0:64]),
		.cby_4__2__chany_top_in(tile_4__2__8_sb_4__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[10]),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__7_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_4__1__chanx_right_out(tile_4__2__7_sb_4__1__chanx_right_out[0:64]),
		.sb_4__1__chany_bottom_out(tile_4__2__7_sb_4__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_4__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__7_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_4__1__chanx_left_out(tile_4__2__7_cbx_4__1__chanx_left_out[0:64]),
		.cby_4__2__chany_top_out(tile_4__2__7_cby_4__2__chany_top_out[0:64]),
		.ccff_tail(tile_4__2__7_ccff_tail));

	tile_4__2_ tile_5__3_ (
		.prog_clk(prog_clk),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_6__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_6__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_6__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_6__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_6__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_6__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__7_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__chanx_right_in(tile_6__2__1_cbx_6__1__chanx_left_out[0:64]),
		.sb_4__1__chany_bottom_in(tile_4__2__7_cby_4__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_16_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_4__1__chanx_left_in(tile_4__2__1_sb_4__1__chanx_right_out[0:64]),
		.cby_4__2__chany_top_in(tile_4__2__9_sb_4__1__chany_bottom_out[0:64]),
		.ccff_head(tile_6__2__1_ccff_tail),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__8_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_4__1__chanx_right_out(tile_4__2__8_sb_4__1__chanx_right_out[0:64]),
		.sb_4__1__chany_bottom_out(tile_4__2__8_sb_4__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_4__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__8_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_4__1__chanx_left_out(tile_4__2__8_cbx_4__1__chanx_left_out[0:64]),
		.cby_4__2__chany_top_out(tile_4__2__8_cby_4__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[13]));

	tile_4__2_ tile_5__4_ (
		.prog_clk(prog_clk),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_6__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_6__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_6__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_6__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_6__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_6__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__8_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__chanx_right_in(tile_6__2__2_cbx_6__1__chanx_left_out[0:64]),
		.sb_4__1__chany_bottom_in(tile_4__2__8_cby_4__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_17_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_4__1__chanx_left_in(tile_4__2__2_sb_4__1__chanx_right_out[0:64]),
		.cby_4__2__chany_top_in(tile_4__2__10_sb_4__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[18]),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__9_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_4__1__chanx_right_out(tile_4__2__9_sb_4__1__chanx_right_out[0:64]),
		.sb_4__1__chany_bottom_out(tile_4__2__9_sb_4__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_4__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__9_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_4__1__chanx_left_out(tile_4__2__9_cbx_4__1__chanx_left_out[0:64]),
		.cby_4__2__chany_top_out(tile_4__2__9_cby_4__2__chany_top_out[0:64]),
		.ccff_tail(tile_4__2__9_ccff_tail));

	tile_4__2_ tile_5__5_ (
		.prog_clk(prog_clk),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_6__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_6__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_6__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_6__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_6__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_6__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__9_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__chanx_right_in(tile_6__2__3_cbx_6__1__chanx_left_out[0:64]),
		.sb_4__1__chany_bottom_in(tile_4__2__9_cby_4__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_18_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_4__1__chanx_left_in(tile_4__2__3_sb_4__1__chanx_right_out[0:64]),
		.cby_4__2__chany_top_in(tile_4__2__11_sb_4__1__chany_bottom_out[0:64]),
		.ccff_head(tile_6__2__3_ccff_tail),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__10_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_4__1__chanx_right_out(tile_4__2__10_sb_4__1__chanx_right_out[0:64]),
		.sb_4__1__chany_bottom_out(tile_4__2__10_sb_4__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_4__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__10_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_4__1__chanx_left_out(tile_4__2__10_cbx_4__1__chanx_left_out[0:64]),
		.cby_4__2__chany_top_out(tile_4__2__10_cby_4__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[21]));

	tile_4__2_ tile_5__6_ (
		.prog_clk(prog_clk),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_6__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_6__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_6__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_6__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_6__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_6__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__10_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__chanx_right_in(tile_6__2__4_cbx_6__1__chanx_left_out[0:64]),
		.sb_4__1__chany_bottom_in(tile_4__2__10_cby_4__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_19_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_4__1__chanx_left_in(tile_4__2__4_sb_4__1__chanx_right_out[0:64]),
		.cby_4__2__chany_top_in(tile_4__2__12_sb_4__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[26]),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__11_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_4__1__chanx_right_out(tile_4__2__11_sb_4__1__chanx_right_out[0:64]),
		.sb_4__1__chany_bottom_out(tile_4__2__11_sb_4__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_4__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__11_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_4__1__chanx_left_out(tile_4__2__11_cbx_4__1__chanx_left_out[0:64]),
		.cby_4__2__chany_top_out(tile_4__2__11_cby_4__2__chany_top_out[0:64]),
		.ccff_tail(tile_4__2__11_ccff_tail));

	tile_4__2_ tile_5__7_ (
		.prog_clk(prog_clk),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_6__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_6__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_6__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_6__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_6__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_6__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__11_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__chanx_right_in(tile_6__2__5_cbx_6__1__chanx_left_out[0:64]),
		.sb_4__1__chany_bottom_in(tile_4__2__11_cby_4__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_20_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_4__1__chanx_left_in(tile_4__2__5_sb_4__1__chanx_right_out[0:64]),
		.cby_4__2__chany_top_in(tile_4__2__13_sb_4__1__chany_bottom_out[0:64]),
		.ccff_head(tile_6__2__5_ccff_tail),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__12_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_4__1__chanx_right_out(tile_4__2__12_sb_4__1__chanx_right_out[0:64]),
		.sb_4__1__chany_bottom_out(tile_4__2__12_sb_4__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_4__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__12_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_4__1__chanx_left_out(tile_4__2__12_cbx_4__1__chanx_left_out[0:64]),
		.cby_4__2__chany_top_out(tile_4__2__12_cby_4__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[29]));

	tile_4__2_ tile_5__8_ (
		.prog_clk(prog_clk),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_6__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_6__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_6__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_6__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_6__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.sb_4__1__right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_6__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_4__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_4__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__12_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_4__1__chanx_right_in(tile_6__2__6_cbx_6__1__chanx_left_out[0:64]),
		.sb_4__1__chany_bottom_in(tile_4__2__12_cby_4__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__9__1_cbx_4__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_5__8__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_4__1__chanx_left_in(tile_4__2__6_sb_4__1__chanx_right_out[0:64]),
		.cby_4__2__chany_top_in(tile_4__9__1_sb_4__8__chany_bottom_out[0:64]),
		.ccff_head(tile_4__2__6_ccff_tail),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_4__2__13_cbx_4__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_4__1__chanx_right_out(tile_4__2__13_sb_4__1__chanx_right_out[0:64]),
		.sb_4__1__chany_bottom_out(tile_4__2__13_sb_4__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_4__2__13_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_4__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_4__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_4__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_4__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_4__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_4__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_4__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_4__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_4__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_4__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_4__2__13_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_4__1__chanx_left_out(tile_4__2__13_cbx_4__1__chanx_left_out[0:64]),
		.cby_4__2__chany_top_out(tile_4__2__13_cby_4__2__chany_top_out[0:64]),
		.ccff_tail(tile_4__2__13_ccff_tail));

	tile_6__1_ tile_6__1_ (
		.prog_clk(prog_clk),
		.sb_6__0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__1_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_6__0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__1_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_6__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__2_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_6__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__2_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_6__0__chanx_right_in(tile_7__1__0_cbx_7__0__chanx_left_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_21_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_6__0__chanx_left_in(tile_4__1__1_sb_4__0__chanx_right_out[0:64]),
		.cby_6__1__chany_top_in(tile_6__2__0_sb_6__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[5]),
		.cbx_6__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_6__1__0_cbx_6__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_6__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_6__1__0_cbx_6__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_6__0__chanx_right_out(tile_6__1__0_sb_6__0__chanx_right_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_6__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_6__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_6__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_6__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_6__1__undriven_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_6__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_6__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_6__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_6__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_6__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_6__1__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_6__0__chanx_left_out(tile_6__1__0_cbx_6__0__chanx_left_out[0:64]),
		.cby_6__1__chany_top_out(tile_6__1__0_cby_6__1__chany_top_out[0:64]),
		.ccff_tail(tile_6__1__0_ccff_tail));

	tile_6__2_ tile_6__2_ (
		.prog_clk(prog_clk),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_6__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_6__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_6__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_6__1__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__1__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_6__1__chanx_right_in(tile_7__2__0_cbx_7__1__chanx_left_out[0:64]),
		.sb_6__1__chany_bottom_in(tile_6__1__0_cby_6__1__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_22_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_6__1__chanx_left_in(tile_4__2__7_sb_4__1__chanx_right_out[0:64]),
		.cby_6__2__chany_top_in(tile_6__2__1_sb_6__1__chany_bottom_out[0:64]),
		.ccff_head(tile_4__2__7_ccff_tail),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_6__2__0_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_6__1__chanx_right_out(tile_6__2__0_sb_6__1__chanx_right_out[0:64]),
		.sb_6__1__chany_bottom_out(tile_6__2__0_sb_6__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_6__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_6__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_6__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_6__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_6__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_6__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_6__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_6__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_6__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_6__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_6__2__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_6__1__chanx_left_out(tile_6__2__0_cbx_6__1__chanx_left_out[0:64]),
		.cby_6__2__chany_top_out(tile_6__2__0_cby_6__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[10]));

	tile_6__2_ tile_6__3_ (
		.prog_clk(prog_clk),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_6__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_6__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_6__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_6__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_6__1__chanx_right_in(tile_7__2__1_cbx_7__1__chanx_left_out[0:64]),
		.sb_6__1__chany_bottom_in(tile_6__2__0_cby_6__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_23_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_6__1__chanx_left_in(tile_4__2__8_sb_4__1__chanx_right_out[0:64]),
		.cby_6__2__chany_top_in(tile_6__2__2_sb_6__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[13]),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_6__2__1_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_6__1__chanx_right_out(tile_6__2__1_sb_6__1__chanx_right_out[0:64]),
		.sb_6__1__chany_bottom_out(tile_6__2__1_sb_6__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_6__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_6__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_6__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_6__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_6__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_6__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_6__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_6__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_6__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_6__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_6__2__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_6__1__chanx_left_out(tile_6__2__1_cbx_6__1__chanx_left_out[0:64]),
		.cby_6__2__chany_top_out(tile_6__2__1_cby_6__2__chany_top_out[0:64]),
		.ccff_tail(tile_6__2__1_ccff_tail));

	tile_6__2_ tile_6__4_ (
		.prog_clk(prog_clk),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_6__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_6__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_6__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_6__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_6__1__chanx_right_in(tile_7__2__2_cbx_7__1__chanx_left_out[0:64]),
		.sb_6__1__chany_bottom_in(tile_6__2__1_cby_6__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_24_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_6__1__chanx_left_in(tile_4__2__9_sb_4__1__chanx_right_out[0:64]),
		.cby_6__2__chany_top_in(tile_6__2__3_sb_6__1__chany_bottom_out[0:64]),
		.ccff_head(tile_4__2__9_ccff_tail),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_6__2__2_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_6__1__chanx_right_out(tile_6__2__2_sb_6__1__chanx_right_out[0:64]),
		.sb_6__1__chany_bottom_out(tile_6__2__2_sb_6__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_6__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_6__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_6__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_6__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_6__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_6__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_6__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_6__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_6__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_6__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_6__2__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_6__1__chanx_left_out(tile_6__2__2_cbx_6__1__chanx_left_out[0:64]),
		.cby_6__2__chany_top_out(tile_6__2__2_cby_6__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[18]));

	tile_6__2_ tile_6__5_ (
		.prog_clk(prog_clk),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_6__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_6__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_6__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_6__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_6__1__chanx_right_in(tile_7__2__3_cbx_7__1__chanx_left_out[0:64]),
		.sb_6__1__chany_bottom_in(tile_6__2__2_cby_6__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_25_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_6__1__chanx_left_in(tile_4__2__10_sb_4__1__chanx_right_out[0:64]),
		.cby_6__2__chany_top_in(tile_6__2__4_sb_6__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[21]),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_6__2__3_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_6__1__chanx_right_out(tile_6__2__3_sb_6__1__chanx_right_out[0:64]),
		.sb_6__1__chany_bottom_out(tile_6__2__3_sb_6__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_6__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_6__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_6__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_6__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_6__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_6__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_6__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_6__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_6__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_6__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_6__2__3_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_6__1__chanx_left_out(tile_6__2__3_cbx_6__1__chanx_left_out[0:64]),
		.cby_6__2__chany_top_out(tile_6__2__3_cby_6__2__chany_top_out[0:64]),
		.ccff_tail(tile_6__2__3_ccff_tail));

	tile_6__2_ tile_6__6_ (
		.prog_clk(prog_clk),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_6__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_6__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_6__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_6__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__3_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_6__1__chanx_right_in(tile_7__2__4_cbx_7__1__chanx_left_out[0:64]),
		.sb_6__1__chany_bottom_in(tile_6__2__3_cby_6__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_26_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_6__1__chanx_left_in(tile_4__2__11_sb_4__1__chanx_right_out[0:64]),
		.cby_6__2__chany_top_in(tile_6__2__5_sb_6__1__chany_bottom_out[0:64]),
		.ccff_head(tile_4__2__11_ccff_tail),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_6__2__4_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_6__1__chanx_right_out(tile_6__2__4_sb_6__1__chanx_right_out[0:64]),
		.sb_6__1__chany_bottom_out(tile_6__2__4_sb_6__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_6__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_6__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_6__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_6__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_6__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_6__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_6__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_6__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_6__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_6__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_6__2__4_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_6__1__chanx_left_out(tile_6__2__4_cbx_6__1__chanx_left_out[0:64]),
		.cby_6__2__chany_top_out(tile_6__2__4_cby_6__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[26]));

	tile_6__2_ tile_6__7_ (
		.prog_clk(prog_clk),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_6__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_6__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_6__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_6__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__4_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_6__1__chanx_right_in(tile_7__2__5_cbx_7__1__chanx_left_out[0:64]),
		.sb_6__1__chany_bottom_in(tile_6__2__4_cby_6__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_27_out),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_6__1__chanx_left_in(tile_4__2__12_sb_4__1__chanx_right_out[0:64]),
		.cby_6__2__chany_top_in(tile_6__2__6_sb_6__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[29]),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_6__2__5_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_6__1__chanx_right_out(tile_6__2__5_sb_6__1__chanx_right_out[0:64]),
		.sb_6__1__chany_bottom_out(tile_6__2__5_sb_6__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_6__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_6__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_6__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_6__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_6__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_6__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_6__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_6__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_6__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_6__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_6__2__5_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_6__1__chanx_left_out(tile_6__2__5_cbx_6__1__chanx_left_out[0:64]),
		.cby_6__2__chany_top_out(tile_6__2__5_cby_6__2__chany_top_out[0:64]),
		.ccff_tail(tile_6__2__5_ccff_tail));

	tile_6__2_ tile_6__8_ (
		.prog_clk(prog_clk),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_6__1__right_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_6__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_6__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_6__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_6__1__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_6__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.sb_6__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__5_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.sb_6__1__chanx_right_in(tile_7__2__6_cbx_7__1__chanx_left_out[0:64]),
		.sb_6__1__chany_bottom_in(tile_6__2__5_cby_6__2__chany_top_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_0_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0_1_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_0_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1_1_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_0_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2_1_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_6__9__0_cbx_6__8__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_(tile_6__8__undriven_grid_clb_left_width_0_height_0_subtile_0__pin_cin_0_),
		.grid_clb_left_width_0_height_0_subtile_0__pin_reset_0_(Reset),
		.grid_clb_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_6__1__chanx_left_in(tile_4__2__13_sb_4__1__chanx_right_out[0:64]),
		.cby_6__2__chany_top_in(tile_6__9__0_sb_6__8__chany_bottom_out[0:64]),
		.ccff_head(tile_4__2__13_ccff_tail),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(tile_6__2__6_cbx_6__1__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.sb_6__1__chanx_right_out(tile_6__2__6_sb_6__1__chanx_right_out[0:64]),
		.sb_6__1__chany_bottom_out(tile_6__2__6_sb_6__1__chany_bottom_out[0:64]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_0_(tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_1_(tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_2_(tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_3_(tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_4_(tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_5_(tile_6__2__6_grid_clb_top_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_6__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_6__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_6__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_6__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_(tile_6__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_(tile_6__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_(tile_6__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_(tile_6__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_(tile_6__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_(tile_6__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_(tile_6__2__6_grid_clb_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.cbx_6__1__chanx_left_out(tile_6__2__6_cbx_6__1__chanx_left_out[0:64]),
		.cby_6__2__chany_top_out(tile_6__2__6_cby_6__2__chany_top_out[0:64]),
		.ccff_tail(tile_6__2__6_ccff_tail));

	tile_7__1_ tile_7__1_ (
		.prog_clk(prog_clk),
		.sb_7__0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__0_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_7__0__right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__0_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_7__0__left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__1_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_7__0__left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__1_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_8__0__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__7_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_8__0__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__7_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_8__0__left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(tile_1__0__0_grid_io_bottom_bottom_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_8__0__left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(tile_1__0__0_grid_io_bottom_bottom_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_7__0__chanx_left_in(tile_6__1__0_sb_6__0__chanx_right_out[0:64]),
		.cby_8__1__chany_top_in(tile_7__2__0_sb_8__1__chany_bottom_out[0:64]),
		.ccff_head(tile_9__1__7_ccff_tail),
		.cbx_7__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__1__0_cbx_7__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_7__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__1__0_cbx_7__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.cbx_8__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__1__0_cbx_8__0__bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.cbx_8__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__1__0_cbx_8__0__bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.cby_8__1__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__1__0_cby_8__1__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_8__1__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__1__0_cby_8__1__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_7__0__chanx_left_out(tile_7__1__0_cbx_7__0__chanx_left_out[0:64]),
		.cby_8__1__chany_top_out(tile_7__1__0_cby_8__1__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[4]));

	tile_7__2_ tile_7__2_ (
		.prog_clk(prog_clk),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__1__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_8__1__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__6_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_8__1__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__6_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_8__1__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__7_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_8__1__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__7_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_8__1__chany_bottom_in(tile_7__1__0_cby_8__1__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_7__1__chanx_left_in(tile_6__2__0_sb_6__1__chanx_right_out[0:64]),
		.cby_8__2__chany_top_in(tile_7__2__1_sb_8__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[11]),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_7__2__0_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__2__0_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__2__0_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_8__1__chany_bottom_out(tile_7__2__0_sb_8__1__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_7__1__chanx_left_out(tile_7__2__0_cbx_7__1__chanx_left_out[0:64]),
		.cby_8__2__chany_top_out(tile_7__2__0_cby_8__2__chany_top_out[0:64]),
		.ccff_tail(tile_7__2__0_ccff_tail));

	tile_7__2_ tile_7__3_ (
		.prog_clk(prog_clk),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__0_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_8__1__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__5_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_8__1__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__5_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_8__1__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__6_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_8__1__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__6_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_8__1__chany_bottom_in(tile_7__2__0_cby_8__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_7__1__chanx_left_in(tile_6__2__1_sb_6__1__chanx_right_out[0:64]),
		.cby_8__2__chany_top_in(tile_7__2__2_sb_8__1__chany_bottom_out[0:64]),
		.ccff_head(tile_9__1__5_ccff_tail),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_7__2__1_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__2__1_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__2__1_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_8__1__chany_bottom_out(tile_7__2__1_sb_8__1__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_7__1__chanx_left_out(tile_7__2__1_cbx_7__1__chanx_left_out[0:64]),
		.cby_8__2__chany_top_out(tile_7__2__1_cby_8__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[12]));

	tile_7__2_ tile_7__4_ (
		.prog_clk(prog_clk),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__1_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_8__1__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__4_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_8__1__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__4_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_8__1__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__5_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_8__1__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__5_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_8__1__chany_bottom_in(tile_7__2__1_cby_8__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_7__1__chanx_left_in(tile_6__2__2_sb_6__1__chanx_right_out[0:64]),
		.cby_8__2__chany_top_in(tile_7__2__3_sb_8__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[19]),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_7__2__2_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__2__2_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__2__2_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_8__1__chany_bottom_out(tile_7__2__2_sb_8__1__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_7__1__chanx_left_out(tile_7__2__2_cbx_7__1__chanx_left_out[0:64]),
		.cby_8__2__chany_top_out(tile_7__2__2_cby_8__2__chany_top_out[0:64]),
		.ccff_tail(tile_7__2__2_ccff_tail));

	tile_7__2_ tile_7__5_ (
		.prog_clk(prog_clk),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__2_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_8__1__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__3_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_8__1__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__3_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_8__1__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__4_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_8__1__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__4_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_8__1__chany_bottom_in(tile_7__2__2_cby_8__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_7__1__chanx_left_in(tile_6__2__3_sb_6__1__chanx_right_out[0:64]),
		.cby_8__2__chany_top_in(tile_7__2__4_sb_8__1__chany_bottom_out[0:64]),
		.ccff_head(tile_9__1__3_ccff_tail),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_7__2__3_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__2__3_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__2__3_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_8__1__chany_bottom_out(tile_7__2__3_sb_8__1__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_7__1__chanx_left_out(tile_7__2__3_cbx_7__1__chanx_left_out[0:64]),
		.cby_8__2__chany_top_out(tile_7__2__3_cby_8__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[20]));

	tile_7__2_ tile_7__6_ (
		.prog_clk(prog_clk),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__3_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_8__1__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__2_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_8__1__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__2_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_8__1__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__3_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_8__1__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__3_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_8__1__chany_bottom_in(tile_7__2__3_cby_8__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_7__1__chanx_left_in(tile_6__2__4_sb_6__1__chanx_right_out[0:64]),
		.cby_8__2__chany_top_in(tile_7__2__5_sb_8__1__chany_bottom_out[0:64]),
		.ccff_head(ccff_head[27]),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_7__2__4_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__2__4_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__2__4_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_8__1__chany_bottom_out(tile_7__2__4_sb_8__1__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_7__1__chanx_left_out(tile_7__2__4_cbx_7__1__chanx_left_out[0:64]),
		.cby_8__2__chany_top_out(tile_7__2__4_cby_8__2__chany_top_out[0:64]),
		.ccff_tail(tile_7__2__4_ccff_tail));

	tile_7__2_ tile_7__7_ (
		.prog_clk(prog_clk),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__4_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_8__1__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__1_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_8__1__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__1_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_8__1__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__2_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_8__1__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__2_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_8__1__chany_bottom_in(tile_7__2__4_cby_8__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_7__1__chanx_left_in(tile_6__2__5_sb_6__1__chanx_right_out[0:64]),
		.cby_8__2__chany_top_in(tile_7__2__6_sb_8__1__chany_bottom_out[0:64]),
		.ccff_head(tile_9__1__1_ccff_tail),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_7__2__5_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__2__5_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__2__5_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_8__1__chany_bottom_out(tile_7__2__5_sb_8__1__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_7__1__chanx_left_out(tile_7__2__5_cbx_7__1__chanx_left_out[0:64]),
		.cby_8__2__chany_top_out(tile_7__2__5_cby_8__2__chany_top_out[0:64]),
		.ccff_tail(ccff_tail[28]));

	tile_7__2_ tile_7__8_ (
		.prog_clk(prog_clk),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.sb_7__1__left_bottom_grid_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__5_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.sb_8__1__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__0_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_8__1__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__0_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_8__1__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(tile_9__1__1_grid_io_right_right_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.sb_8__1__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(tile_9__1__1_grid_io_right_right_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.sb_8__1__chany_bottom_in(tile_7__2__5_cby_8__2__chany_top_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_7__9__0_cbx_7__8__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.grid_memory_left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.cbx_7__1__chanx_left_in(tile_6__2__6_sb_6__1__chanx_right_out[0:64]),
		.cby_8__2__chany_top_in(tile_8__9__0_sb_8__8__chany_bottom_out[0:64]),
		.ccff_head(tile_6__2__6_ccff_tail),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_(tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_0_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_(tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_1_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_(tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_2_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_(tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_3_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_(tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_4_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_(tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_5_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_(tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_6_),
		.cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_(tile_7__2__6_cbx_7__1__bottom_grid_top_width_0_height_0_subtile_0__pin_d_in_7_),
		.cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(tile_7__2__6_cby_8__2__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(tile_7__2__6_cby_8__2__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.sb_8__1__chany_bottom_out(tile_7__2__6_sb_8__1__chany_bottom_out[0:64]),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_0_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_1_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_2_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_3_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_4_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_5_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_6_),
		.grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_(tile_7__2__6_grid_memory_top_width_0_height_0_subtile_0__pin_d_out_7_),
		.cbx_7__1__chanx_left_out(tile_7__2__6_cbx_7__1__chanx_left_out[0:64]),
		.cby_8__2__chany_top_out(tile_7__2__6_cby_8__2__chany_top_out[0:64]),
		.ccff_tail(tile_7__2__6_ccff_tail));

	direct_interc direct_interc_0_ (
		.in(tile_1__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_0_out));

	direct_interc direct_interc_1_ (
		.in(tile_1__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_1_out));

	direct_interc direct_interc_2_ (
		.in(tile_1__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_2_out));

	direct_interc direct_interc_3_ (
		.in(tile_1__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_3_out));

	direct_interc direct_interc_4_ (
		.in(tile_1__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_4_out));

	direct_interc direct_interc_5_ (
		.in(tile_1__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_5_out));

	direct_interc direct_interc_6_ (
		.in(tile_1__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_6_out));

	direct_interc direct_interc_7_ (
		.in(tile_4__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_7_out));

	direct_interc direct_interc_8_ (
		.in(tile_4__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_8_out));

	direct_interc direct_interc_9_ (
		.in(tile_4__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_9_out));

	direct_interc direct_interc_10_ (
		.in(tile_4__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_10_out));

	direct_interc direct_interc_11_ (
		.in(tile_4__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_11_out));

	direct_interc direct_interc_12_ (
		.in(tile_4__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_12_out));

	direct_interc direct_interc_13_ (
		.in(tile_4__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_13_out));

	direct_interc direct_interc_14_ (
		.in(tile_4__2__7_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_14_out));

	direct_interc direct_interc_15_ (
		.in(tile_4__2__8_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_15_out));

	direct_interc direct_interc_16_ (
		.in(tile_4__2__9_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_16_out));

	direct_interc direct_interc_17_ (
		.in(tile_4__2__10_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_17_out));

	direct_interc direct_interc_18_ (
		.in(tile_4__2__11_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_18_out));

	direct_interc direct_interc_19_ (
		.in(tile_4__2__12_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_19_out));

	direct_interc direct_interc_20_ (
		.in(tile_4__2__13_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_20_out));

	direct_interc direct_interc_21_ (
		.in(tile_6__2__0_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_21_out));

	direct_interc direct_interc_22_ (
		.in(tile_6__2__1_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_22_out));

	direct_interc direct_interc_23_ (
		.in(tile_6__2__2_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_23_out));

	direct_interc direct_interc_24_ (
		.in(tile_6__2__3_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_24_out));

	direct_interc direct_interc_25_ (
		.in(tile_6__2__4_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_25_out));

	direct_interc direct_interc_26_ (
		.in(tile_6__2__5_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_26_out));

	direct_interc direct_interc_27_ (
		.in(tile_6__2__6_grid_clb_right_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_27_out));

endmodule
// ----- END Verilog module for fpga_top -----

//----- Default net type -----
`default_nettype wire




