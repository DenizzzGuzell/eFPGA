//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Tile Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed Aug 14 09:11:37 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype wire

// ----- Verilog module for tile_17__10_ -----
module tile_17__10_(prog_clk,
                    sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
                    sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_,
                    sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                    sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_,
                    sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
                    sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_,
                    sb_17__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_,
                    sb_17__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_,
                    sb_17__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_,
                    sb_17__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_,
                    sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
                    sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_,
                    sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                    sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_,
                    sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
                    sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_,
                    sb_18__9__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
                    sb_18__9__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
                    sb_18__9__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
                    sb_18__9__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
                    sb_18__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_,
                    sb_18__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_,
                    sb_18__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_,
                    sb_18__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_,
                    sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
                    sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_,
                    sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                    sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_,
                    sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
                    sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_,
                    sb_17__9__chany_bottom_in,
                    sb_18__9__chany_bottom_in,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_,
                    grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_,
                    cbx_17__9__chanx_left_in,
                    cby_18__10__chany_top_in,
                    ccff_head,
                    cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_,
                    cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_,
                    cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_,
                    cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_,
                    cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_,
                    cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_,
                    cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_,
                    cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_,
                    cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_,
                    cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_,
                    cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_,
                    cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_,
                    cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_,
                    cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_,
                    cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_,
                    cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_,
                    cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_,
                    cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_,
                    cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_,
                    cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_,
                    cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_,
                    cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_,
                    cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_,
                    cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_,
                    cby_18__10__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_,
                    cby_18__10__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_,
                    sb_17__9__chany_bottom_out,
                    sb_18__9__chany_bottom_out,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_,
                    grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_,
                    cbx_17__9__chanx_left_out,
                    cby_18__10__chany_top_out,
                    ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
//----- INPUT PORTS -----
input [0:0] sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_;
//----- INPUT PORTS -----
input [0:0] sb_17__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
//----- INPUT PORTS -----
input [0:0] sb_17__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
//----- INPUT PORTS -----
input [0:0] sb_17__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
//----- INPUT PORTS -----
input [0:0] sb_17__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
//----- INPUT PORTS -----
input [0:0] sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
//----- INPUT PORTS -----
input [0:0] sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_;
//----- INPUT PORTS -----
input [0:0] sb_18__9__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] sb_18__9__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] sb_18__9__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] sb_18__9__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] sb_18__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
//----- INPUT PORTS -----
input [0:0] sb_18__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
//----- INPUT PORTS -----
input [0:0] sb_18__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
//----- INPUT PORTS -----
input [0:0] sb_18__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
//----- INPUT PORTS -----
input [0:0] sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
//----- INPUT PORTS -----
input [0:0] sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_;
//----- INPUT PORTS -----
input [0:64] sb_17__9__chany_bottom_in;
//----- INPUT PORTS -----
input [0:64] sb_18__9__chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_;
//----- INPUT PORTS -----
input [0:0] grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_;
//----- INPUT PORTS -----
input [0:64] cbx_17__9__chanx_left_in;
//----- INPUT PORTS -----
input [0:64] cby_18__10__chany_top_in;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_;
//----- OUTPUT PORTS -----
output [0:0] cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_;
//----- OUTPUT PORTS -----
output [0:0] cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_;
//----- OUTPUT PORTS -----
output [0:0] cby_18__10__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
//----- OUTPUT PORTS -----
output [0:0] cby_18__10__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
//----- OUTPUT PORTS -----
output [0:64] sb_17__9__chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:64] sb_18__9__chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_;
//----- OUTPUT PORTS -----
output [0:0] grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_;
//----- OUTPUT PORTS -----
output [0:64] cbx_17__9__chanx_left_out;
//----- OUTPUT PORTS -----
output [0:64] cby_18__10__chany_top_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:0] cbx_1__9__0_ccff_tail;
wire [0:64] cbx_1__9__0_chanx_right_out;
wire [0:0] cbx_1__9__1_ccff_tail;
wire [0:64] cbx_1__9__1_chanx_left_out;
wire [0:64] cbx_1__9__1_chanx_right_out;
wire [0:0] cby_18__5__0_ccff_tail;
wire [0:64] cby_18__5__0_chany_bottom_out;
wire [0:64] sb_18__4__0_chanx_left_out;
wire [0:64] sb_18__4__0_chany_top_out;
wire [0:0] sb_1__9__0_ccff_tail;
wire [0:64] sb_1__9__0_chanx_left_out;
wire [0:64] sb_1__9__0_chanx_right_out;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	grid_mult_18 grid_mult_18_17__10_ (
		.top_width_0_height_0_subtile_0__pin_sign_0_(grid_mult_18_top_width_0_height_0_subtile_0__pin_sign_0_),
		.top_width_0_height_0_subtile_0__pin_a_0_(grid_mult_18_top_width_0_height_0_subtile_0__pin_a_0_),
		.top_width_0_height_0_subtile_0__pin_a_1_(grid_mult_18_top_width_0_height_0_subtile_0__pin_a_1_),
		.top_width_0_height_0_subtile_0__pin_a_2_(grid_mult_18_top_width_0_height_0_subtile_0__pin_a_2_),
		.top_width_0_height_0_subtile_0__pin_a_3_(grid_mult_18_top_width_0_height_0_subtile_0__pin_a_3_),
		.top_width_0_height_0_subtile_0__pin_a_4_(grid_mult_18_top_width_0_height_0_subtile_0__pin_a_4_),
		.top_width_0_height_0_subtile_0__pin_a_5_(grid_mult_18_top_width_0_height_0_subtile_0__pin_a_5_),
		.top_width_0_height_0_subtile_0__pin_a_6_(grid_mult_18_top_width_0_height_0_subtile_0__pin_a_6_),
		.top_width_0_height_0_subtile_0__pin_a_7_(grid_mult_18_top_width_0_height_0_subtile_0__pin_a_7_),
		.top_width_0_height_0_subtile_0__pin_a_8_(grid_mult_18_top_width_0_height_0_subtile_0__pin_a_8_),
		.top_width_0_height_0_subtile_0__pin_a_9_(grid_mult_18_top_width_0_height_0_subtile_0__pin_a_9_),
		.top_width_0_height_0_subtile_0__pin_a_10_(grid_mult_18_top_width_0_height_0_subtile_0__pin_a_10_),
		.top_width_0_height_0_subtile_0__pin_a_11_(grid_mult_18_top_width_0_height_0_subtile_0__pin_a_11_),
		.top_width_0_height_0_subtile_0__pin_a_12_(grid_mult_18_top_width_0_height_0_subtile_0__pin_a_12_),
		.top_width_0_height_0_subtile_0__pin_a_13_(grid_mult_18_top_width_0_height_0_subtile_0__pin_a_13_),
		.top_width_0_height_0_subtile_0__pin_a_14_(grid_mult_18_top_width_0_height_0_subtile_0__pin_a_14_),
		.top_width_0_height_0_subtile_0__pin_a_15_(grid_mult_18_top_width_0_height_0_subtile_0__pin_a_15_),
		.top_width_0_height_0_subtile_0__pin_a_16_(grid_mult_18_top_width_0_height_0_subtile_0__pin_a_16_),
		.top_width_0_height_0_subtile_0__pin_a_17_(grid_mult_18_top_width_0_height_0_subtile_0__pin_a_17_),
		.top_width_0_height_0_subtile_0__pin_a_18_(grid_mult_18_top_width_0_height_0_subtile_0__pin_a_18_),
		.top_width_0_height_0_subtile_0__pin_b_0_(grid_mult_18_top_width_0_height_0_subtile_0__pin_b_0_),
		.top_width_0_height_0_subtile_0__pin_b_1_(grid_mult_18_top_width_0_height_0_subtile_0__pin_b_1_),
		.top_width_0_height_0_subtile_0__pin_b_2_(grid_mult_18_top_width_0_height_0_subtile_0__pin_b_2_),
		.top_width_0_height_0_subtile_0__pin_b_3_(grid_mult_18_top_width_0_height_0_subtile_0__pin_b_3_),
		.top_width_0_height_0_subtile_0__pin_b_4_(grid_mult_18_top_width_0_height_0_subtile_0__pin_b_4_),
		.top_width_0_height_0_subtile_0__pin_b_5_(grid_mult_18_top_width_0_height_0_subtile_0__pin_b_5_),
		.top_width_0_height_0_subtile_0__pin_b_6_(grid_mult_18_top_width_0_height_0_subtile_0__pin_b_6_),
		.top_width_0_height_0_subtile_0__pin_b_7_(grid_mult_18_top_width_0_height_0_subtile_0__pin_b_7_),
		.top_width_0_height_0_subtile_0__pin_b_8_(grid_mult_18_top_width_0_height_0_subtile_0__pin_b_8_),
		.top_width_0_height_0_subtile_0__pin_b_9_(grid_mult_18_top_width_0_height_0_subtile_0__pin_b_9_),
		.top_width_0_height_0_subtile_0__pin_b_10_(grid_mult_18_top_width_0_height_0_subtile_0__pin_b_10_),
		.top_width_0_height_0_subtile_0__pin_b_11_(grid_mult_18_top_width_0_height_0_subtile_0__pin_b_11_),
		.top_width_0_height_0_subtile_0__pin_b_12_(grid_mult_18_top_width_0_height_0_subtile_0__pin_b_12_),
		.top_width_0_height_0_subtile_0__pin_b_13_(grid_mult_18_top_width_0_height_0_subtile_0__pin_b_13_),
		.top_width_0_height_0_subtile_0__pin_b_14_(grid_mult_18_top_width_0_height_0_subtile_0__pin_b_14_),
		.top_width_0_height_0_subtile_0__pin_b_15_(grid_mult_18_top_width_0_height_0_subtile_0__pin_b_15_),
		.top_width_0_height_0_subtile_0__pin_b_16_(grid_mult_18_top_width_0_height_0_subtile_0__pin_b_16_),
		.top_width_0_height_0_subtile_0__pin_b_17_(grid_mult_18_top_width_0_height_0_subtile_0__pin_b_17_),
		.top_width_0_height_0_subtile_0__pin_b_18_(grid_mult_18_top_width_0_height_0_subtile_0__pin_b_18_),
		.bottom_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.bottom_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.bottom_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.bottom_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.bottom_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.bottom_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.bottom_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.bottom_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.bottom_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.bottom_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.bottom_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.bottom_width_0_height_0_subtile_0__pin_out_12_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.bottom_width_0_height_0_subtile_0__pin_out_13_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.bottom_width_0_height_0_subtile_0__pin_out_14_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.bottom_width_0_height_0_subtile_0__pin_out_15_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.bottom_width_0_height_0_subtile_0__pin_out_16_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.bottom_width_0_height_0_subtile_0__pin_out_17_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.bottom_width_0_height_0_subtile_0__pin_out_18_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.bottom_width_0_height_0_subtile_0__pin_out_19_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.bottom_width_0_height_0_subtile_0__pin_out_20_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.bottom_width_0_height_0_subtile_0__pin_out_21_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.bottom_width_0_height_0_subtile_0__pin_out_22_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.bottom_width_0_height_0_subtile_0__pin_out_23_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.bottom_width_0_height_0_subtile_0__pin_out_24_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.bottom_width_0_height_0_subtile_0__pin_out_25_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.bottom_width_0_height_0_subtile_0__pin_out_26_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.bottom_width_0_height_0_subtile_0__pin_out_27_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.bottom_width_0_height_0_subtile_0__pin_out_28_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.bottom_width_0_height_0_subtile_0__pin_out_29_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.bottom_width_0_height_0_subtile_0__pin_out_30_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.bottom_width_0_height_0_subtile_0__pin_out_31_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.bottom_width_0_height_0_subtile_0__pin_out_32_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.bottom_width_0_height_0_subtile_0__pin_out_33_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.bottom_width_0_height_0_subtile_0__pin_out_34_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.bottom_width_0_height_0_subtile_0__pin_out_35_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.bottom_width_0_height_0_subtile_0__pin_out_36_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.bottom_width_0_height_0_subtile_0__pin_out_37_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_));

	cbx_1__9_ cbx_17__9_ (
		.prog_clk(prog_clk),
		.chanx_left_in(cbx_17__9__chanx_left_in[0:64]),
		.chanx_right_in(sb_1__9__0_chanx_left_out[0:64]),
		.ccff_head(ccff_head),
		.chanx_left_out(cbx_17__9__chanx_left_out[0:64]),
		.chanx_right_out(cbx_1__9__0_chanx_right_out[0:64]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_17__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.ccff_tail(cbx_1__9__0_ccff_tail));

	cbx_1__9_ cbx_18__9_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__9__0_chanx_right_out[0:64]),
		.chanx_right_in(sb_18__4__0_chanx_left_out[0:64]),
		.ccff_head(cbx_1__9__0_ccff_tail),
		.chanx_left_out(cbx_1__9__1_chanx_left_out[0:64]),
		.chanx_right_out(cbx_1__9__1_chanx_right_out[0:64]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_18__9__bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.ccff_tail(cbx_1__9__1_ccff_tail));

	cby_18__5_ cby_18__10_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_18__4__0_chany_top_out[0:64]),
		.chany_top_in(cby_18__10__chany_top_in[0:64]),
		.ccff_head(cbx_1__9__1_ccff_tail),
		.chany_bottom_out(cby_18__5__0_chany_bottom_out[0:64]),
		.chany_top_out(cby_18__10__chany_top_out[0:64]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_18__10__right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_18__10__right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_tail(cby_18__5__0_ccff_tail));

	sb_1__9_ sb_17__9_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__9__1_chanx_left_out[0:64]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(sb_17__9__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_),
		.chany_bottom_in(sb_17__9__chany_bottom_in[0:64]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_17__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_17__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_17__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_17__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__9__0_chanx_right_out[0:64]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_0_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_1_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_2_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_3_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_3_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_4_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_5_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_6_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_7_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_7_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_8_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_9_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_9_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_10_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_11_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_12_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_13_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_14_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_15_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_16_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_17_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_18_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_19_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_19_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_20_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_21_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_21_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_22_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_22_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_23_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_23_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_24_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_25_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_25_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_26_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_26_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_27_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_27_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_28_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_29_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_29_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_30_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_30_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_31_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_31_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_32_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_33_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_33_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_34_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_34_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_35_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_35_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_36_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_36_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_out_37_(grid_mult_18_bottom_width_0_height_0_subtile_0__pin_out_37_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(sb_17__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_),
		.ccff_head(cby_18__5__0_ccff_tail),
		.chanx_right_out(sb_1__9__0_chanx_right_out[0:64]),
		.chany_bottom_out(sb_17__9__chany_bottom_out[0:64]),
		.chanx_left_out(sb_1__9__0_chanx_left_out[0:64]),
		.ccff_tail(sb_1__9__0_ccff_tail));

	sb_18__4_ sb_18__9_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_18__5__0_chany_bottom_out[0:64]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(sb_18__9__top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(sb_18__9__top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.chany_bottom_in(sb_18__9__chany_bottom_in[0:64]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(sb_18__9__bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(sb_18__9__bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(sb_18__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(sb_18__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(sb_18__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(sb_18__9__bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__9__1_chanx_right_out[0:64]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(sb_18__9__left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_),
		.ccff_head(sb_1__9__0_ccff_tail),
		.chany_top_out(sb_18__4__0_chany_top_out[0:64]),
		.chany_bottom_out(sb_18__9__chany_bottom_out[0:64]),
		.chanx_left_out(sb_18__4__0_chanx_left_out[0:64]),
		.ccff_tail(ccff_tail));

endmodule
// ----- END Verilog module for tile_17__10_ -----

//----- Default net type -----
`default_nettype wire




